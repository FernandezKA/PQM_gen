`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HLBNbspr1A6MAkHQZ9S/syyaXtTVSpkUPj3Wv56LJ6bW6gIzy/56hn7ujs90pFKi6IIk8WLUcAoS
ElGYwvfIrw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
plDDdrKIGUtnra1V+sb5AwOdsrrrHRGchCUGLwrSkI634d818BALn4az/DNSrYPOpdgleXNN3mtS
IKNAXLl9g0B3exvefyuuBenlzYWQXw/8a6ri62ZYhXJfglShAnMwXLb6OMrTffhDBQm15CyqyFei
Rs/au6WGeFoyjM7+fRQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uH+TDuLmzjZd6JKH8ZX4HxGrdBQMKQNF3VaxBr77u09ayo5auQgQmkE8ztTHgo3NMKvY1Z5N+k2W
TRx6wnJo1FmglDEL8XMyLFS8lFjrLeRume7tsdlElfV3kClZjeln8yNgp+Ea3yrlwU2iY477JcoV
J1Iqatzps8xUkTED6cd2SvTYixcPh2wN4D6ojeV9y5IAE+UKQhK3Tn9siQz7swttok5bmLMwzJGo
hKNuakPLTr/MjqCk9A0p/Y4eOCRBrPnvnyqStXpXG8/FUs2LAP+ATQqKLtX9/0/vAFF5qyImKgeE
PVph2EWhSV/Y4tySDMGiziFygukIX+yTp2iGIw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pST7JUFjt9DdbRgc6XMKfp3axHuj4lhmozNUwnyXcVHF+7ATC+DiBF0veEesOZVo+CJaLgEz1SMx
SIeHTZxFjwbr+HrZr3LQknoCL4H2aH7a/+bX22kHT0LxId9UUGkJtuDWVcOhnQxPP3jMdUNq8l99
Ps/y57k6/OrQL9Aa2lIJyGw0rcf31lmaxc6dUlUjVyUwcs8xMAJk3HHtPg4cHzgD9R6LiUR50HB1
ER1ac866L47Fd6sq/Z6sH8WhZtzSlIcyoQWgIFPwtlkKRO/8D5sQ59jLsMa3PUDSelyx5SD+dP0l
nTuDfWpuPSPpItwDH2Q3uYaHS+VU78Dlc3BCrw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YOsQoiX9zSlyfqYxcjGeqz0g/ldv0Zt5FhTqLzdJlgSBH7iwmB8o4Uuxetign7SxzkY+B8IZzNeU
RHfiuwUs+bvDUsJ0s0uSkHfDxGWtzGmOa4ufXS/n0KwEmXJwCmC5s9n0k7UooN0YehoJZ0n2yetb
YylWpoY2NIFF3zrRe9M5fHY6GzDpyHscckrZ4j6coDPoDMEZ4ysK/zXq/91N6IS4ewq1AH3gLa1W
AaxsFJJJCN97KCvky9XfsviK67rHQl0X/9mUmngK0zWrkc8mhIvO/6Le0p4oZwNB/vibZiM/4bPK
BIl9KSo8sEjrbxjr1zUhbGobh2oY90aMFzQmmw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NjCrsxSSgpdJH3xYHdA7jLx598d3jbp0pWnZqMrsEpcm5NoUyOuqQzjnve6v6VnElFWUKuYOm3UB
HUAaCdUqXuXzLtQsCmlGAqlQfsfvprbF9G2t/7Fbi0gZkyyZPTrPH90LOmxYZ2OgDUtthG0pitmv
lxpEV4TFo8smCK8DpY8=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aiMp8Dd5FA+Xh1Vdhf9zMYN/xUTNWlpIcZEBPmzHIGENJ5ofFFhuFckBrYuzH7b2L1DA6oMz6yAW
KDpBkdp/+MCQFbQ2+PFeQHK3C/gl6Mo4shK+YEVg0W9m7ZLrAdyRibP0lv8KxkzDy9ylCI3/E8lx
QVd1bxNhyaYxpXdFXYVwIHQRIeDdIXty4fYHmqHLYuQ04nOmoxqQTBfMKyvIr2nBIIpyMeBAwjq1
a3alou22cPso8teQYrFGTy/WvrwKlwa+0ZFcJ7p+XqY0KqO5G+kFSd0b9UDgx+8YJzyCFjfpp3ds
GeDdbwIeaUATqhNVY4a1suuOMXzz79u7KGdxQg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 96624)
`protect data_block
ijTIFTnqWGCJMMbb3vC/TbrNagFahSdGNyk8xOlEtFgY/RXZaJI7wiy6gGzpOlOUfGtolsCbe6Nz
NijGy7CZ1zHdCfZem6Gj6uuZ5yzA4MyXfiPEwYhD1QKTVmJiFGjEEMvRc+qX1BTcrLYgv5joEa9T
ZAqbgtR3K1ToMAsQY58upLYRkUmTKDvCw5Xy7fCFcnLztSlSk1FMLh3C14J4o3jXajnbVPE8aIyT
8J+NMmk7xx6oqYUXEuLUxqe2zn7aUPCvR6VjJIVxqHwEW3zikoHb1DwUVnZLhR8nanINiSY9dGRL
CyDzyqqpLs1oiYOBK3Lay10gKYfCv4Ope0eYyzpoxMbBJ13y21CXskhs7RpI2iy1TxNIQAld5jj/
bXHjPzJ6uR62wfsQQdLoGJRyhv5I5AhiLD/7KskCKYyX/7j+lxYuDInw3Su/IAUU+i2SbgSUSucg
zvsfbS9n32fTRolWBK7sizZnhDmFZgu4vyV88ZilsEQL7l2ux+OEz/cEOLdRLbdu/og8r08WSYg3
RfnZEaTCxBYzsafO+OENViHsJHYAlkRuGei0BG4LeRjksFQDX51xBm0T+j8t+CHKCpHEf85pvdzc
u6nug9Rkm0nAqyO/POQbY4ttaF+TP5ZHAaRf0n7hVdZ2u4bDv4ROdZel7npdsvXjbgQ9fnkTWxRJ
m40hzn50NiOL03fOI3mfX6lfvjSN4eZGY0fdYIUiNJQn4sMz1TlLyDVyv4iYpfSgq8CPeHaFbJeU
ZzvJRY/Edy0Nbv5GQLYfBPSkKqN3UJgS/rNP5dldWPWHvxmj1xL0BVtIys0I7r/GbyWnLfE+BVex
mzEERTXtearLwP4P/ysh2pt5aw7Fq6Fjxy1zH8NsyzkMgBGxQjBjvaXg20E3fR7cWdPY9th4+oMD
qGCAScfc5Z3La3my683l13cwdf1D0C9N0fGlZvgGpuPe49OMvsENI2k+5vyZGR69gg1dbeZ7YB2l
lq7L6rXZ3y9kqKavCEU8KBmX/PsIKgN3VFQmd8cU32dDTYvkYAYLxnmrH6v1mR768iw5jR+A8fUi
XNYRWQjfSYiW7na8laYUcp2NA2hK2CoiregKjczfgBSlwmX2ATUFAVCbbI32SabMTbMjseN+fkx9
q1QV8rPtCwVo/KR3ramJODULsr6dp62a2So6WdZ6jZaV/jSzH6ZDh4w0jRtw2hzbjvSwg+JVsKCK
2/Oj1yBxNFrbUcAhswdF1AD56IU0Z+IeAZKi/JjcRnQy1P7uraXZsO6Rz4ao+hVKm8Tm8pYq1KsK
OtIaOto9W+OgXmP6iImt0oiXZVppTBJFRNmoRUnxMtjMj9w0iC5b6wxbEZoAFs08j+HScLsWPSHo
dWecBX0zmKBmTy6pPgMXd/NhzIeIQnKpiW2LaPEt8DVUNuE35nkKZaihu5MZxFowhdfZ90S2FI3U
Dw4QVlBhxlBhrH8io7KEVr68Oy1dRMfOd2rtr6BZ669m7eO592VHS/Pcxtjb2cHHv6/t20MUG38l
tgn0y/sj85Gzi8sV7r1mYEiG1yjJl4p+k262AkVTYh6ehMUGoJIolBULTBbk3cEZ28tcRyYStmMm
/G9TLvbz0HU4Lh0Qpng4EXEqUx+ylkLIJ5kw+yAAO4JSVgCsWf4zksxUlX5ez6VK8DLQxk52lG76
EbH8+UvSEpQoZVwp8cCvwIliZl1sf4d4l1Rl4pRL45ht+arX2iiWOs/BqyLNSe8CMIPlkDB+wjfa
jH9oPd9QmUrCokVO1eQYCv3SmW2sLUuZDFP8pANnEj1yZ2T+dXX17MEsHUAkVaHbdBzjMU/XtoaI
SiICgq8Y2XN5IQcpnl5rLjjq4czBDUTH7KE4KwzoRvitOfZJEkAd3aI6IfYDG8kzn+85yFemcH2c
i748iPUKHi3qLBe92THESbDyicD/CsvkR36AYgrQBtDuktg7zJyiPuKHOJfPvAvRxJxdT6hoY8As
Zx2844jXJSf4UXfrdIhMzg7d3cgsShovxzTjxhwazWQ3cmkOUWUM8T8c+AvVn94ZqDa5XRLopDB6
K7vb4h2nFLFu8qYHPs0BWGMMo9xHlskQWzchzDfJIUJ6bgYFjTFvHxx3RvvR+7ybrToYMNTRuoKV
tsaSgadL5S+sNsiWppzTEMBcBMC2xlQeMlQWK6OrIdqoV3IXsejc0rO0SxsYEfXWtwDk78CHlp4I
OMmLO3qAxyvD8SVkG9drPqIy0ZeST+IJN4iEvy0JzrvCi9shI/e2q3D1ej4r82zKwpY1NaC+2d+g
ucCj//2jPTzYLjah2PT8j0q+wTwbQ5n6lrdu6yCydo7gjvaJRJU9M9m1JtPz5/TjkgN/7fgCCEem
tsSX3NLaOWSwXL3zi5/l6vttaGD9yWiQxPABdudPlB8ItUH/lGWqjQbmrC8d0EAOEehL0qW8GaQF
XuVkatpxB+pq5/tDpCNDXjWxW2ednu7yI/19Eik+7hfybD9oz/lFotWSkbwLNbSmlmkwJ2xCWZu6
PRSwzuPJRNiRHs79dga+4oKSnEmfvXRaSQ6eqdNn7oI+XUXunRHSx2x81vk9GzVNjZjWbMTAx6wk
B7dTCl/1YnDOxkHPcGW79KqI1GKgACndo2HwEA3DAzbZUBSBKOnm9yL2PkSlDgaKYrPOMYtLwYT0
yByY/PVLPVy77XDoZZEc40cAujAP/ZTuKot5nDvVuml7HJK6w7CcxyLzB/6LKu1SA3tY80Faoqo1
9TQJYaKTtuVUEhMkdYi8wS5o/qgPbNx5yTY8pSsN/spBwG2mlDz5w9mqtMqHCMHwO2/YKqVskE1+
oVosbNdyVHPs89F49YPGg+rtDLYBJn25yn4Q1C1Tok6wOaVc2IhuUE9b2GJL48QLrdA9zl+OS2Ar
md6cd2+Aqe5nP+Njrm7IICd8qn6hyagQtfmg467OzfOTCMbBPgcq/oSrCSS1oTEQDr4MW4gju6mc
h768WpQDt8qxgpzmQTokCV8k0XWBHfVw6fN5XUvfgS8MnvukGV7WZQ6Y/gJQ9MreuikqOmslB/kk
JCLH6hZrrThoxUuta4k1vkusGqBHuycFg5oeYJjDHHmGJKBb7AAO/gNCLliYLhNlsh+bZGSHqjAw
WpqivXIMhPt/6BERm3tveQi6v8P2Ld4CmeE3XCCch0GCbLtd5+OY0yqhnmqxMzZpvicK+WejostF
n/TJWfZrAHbB4ykbPW48rpoIk6WQdzx8fYEh/fCRVd7XgD1YwvNhxYIplrfNDtcebL0z5R0Kq2jt
IokBtrLgjo5SfQTZXYa6svlPG30dxFCgFO60JUD8w7Hof17iKrIdSuz3Vdp/nCUGgz8Vl0OeLbwY
ojhAeL9G6vhurkbPJ6K5R/0GlnRY69CvMRYag99TDLf3kPav/DOHOg0+KlGFOIiHkHoOcCDAmQ6M
5KU4S63b5/QIAtfkj8WKzauZ2F3dtIBhpPOp8WziXqc9XtvrLS1V9cvp6IQdAtgstZ5g3FjI7vxE
OTr/V5pyixRFWBZnLNN7ZQBjjzWDWAKbsNLfe5uV2/JdbJoibEB1hIaW7G5xtsFa01/tgkT6LS+U
kVezsw3nVibwD9cfRWcMqIrRCwJp6a2Qy6P6iFO+1hvbMNYbIaDcWiZZpE1KiMNwsoiJxskmxkHd
XVmPxo7KR3anvAKI1yq7ye5UYPtiEx161jmK7gpCrG6RgowgZDMAcH+Jn9BjhHeKtdp1CSzvU1I7
NXffmVDWnAdkF9o5W7Lo9yooCAIhk4p/hEmxe0CF2/vwEJLtkBmSItZYeXAFQrx/LtxsF71Ux806
QhiovyDRAbqnxjM2IT5BjIoXriOgSX1OpSedAb/VXhno0gPkwbjiI4iyqGj57L6Z8hs8pWoyHQdB
C1y9T+walO0Du4tvya4rl3OvOLrv6N8kpx5529mZMIVidHbdhxLXSUnh8aquPvIZFCML4q+IVo1q
U6VBhQMIE9aH5H5uJIRML+Ji4miLGRbPWyMDeWVnwVvSF5afUqNIPal/+ugcsj2CyyFeuJjSbxus
j8a8LYq/l4FZfQm3ttzVqIjQnr8V40AWhmh9JDAo+7WVO0CBtimgz/8ylaxeHJMOOdYT/lFq01fz
8romKkOZ8RM09kDbROZt6igI/FuupF2iSG6bU3qEAvAHR7gPgFEEP8Q3fXllPrBbzJHkmoROnbUC
1wRwPfHy1gfEqYJ4FJqPPgcoXo/0NqnHNDnNi70l/nBW0uiLQoVZp5fyyNHea+1EiMxlZp88QsvJ
TK3z+hCbQWqHec4UxQU/nGNbTmERG1BproptbOnIXL53AhzXE2dmTSDQr5P4YVctJ0CHQBLBCHeo
9yifacedEpiyoSomar+PJhYOu3hknev1PcD7USdLTwVAhHAp9mghnyGSNf3EMc72KjPLe1FdjuDR
Ca1djXXUmEeXb5IpRrCNahH+eYWacGoAF9QaxmPVYzYizrwt5jTIIgL2vneL5Ux9DJC35yW7/Obd
TbgjfhTwBdeInWIoKN96+SbLU91idEcfLnOIwlSs6A1RRDNdn2uDFsCGeIANTuNgu4sFLL/DS/F/
hDJwrPXm0ePdNhV+YHNhIEzAFsUn5eceKLWQP5Lyy3mA5LlcHANoreHus58NkB7sxvL3tv63fGGO
SsEXAAh7fBIQXSgETO02N5gsMet9seimsgE/Fe873cdOnJLMRYaBu9NzyiTXjdqKN8bcUET+M0pe
XU1gIaAjlRhyFlQ7pyRmNIRXAL/U/kbx7lW6FWOyAXDQdzlx+UuA3OG4ZDJhofuRYcvcVrpRVQ/1
yYhQVGhHeDXHT/CfoxS67WENReDmraj4IuoaB9MtjO+ijvvDK17x96C0b/MlxZO54EloOzg5xJ4v
T00k462u4gspZZukGPlTCD0I8NBs4PvynMN3IFHiHypSbHiSQiNR1mXuFx5Wjh9EMgXf0pHHH265
g8tl2aYuk8rRnXkbFMZCf1nSEZ47s8PnYZgru8a5fiuhMGpRCVIqGf758UMMMIkXsr0ri7lkr5R1
0HsNUmlBF02dCQq4QLNfYR/WFIYOykAs+S4ofAsPLn0PhXqR+OYhRETONzqhJpImJ5c0K2H3XJjA
WuKNg6yhO0ScUmDMCt6UQPd37zlBWG+baRFFuM0Ih6iUbmEKhQZh3v1lDWueDnWEJr4I72T7gDy2
rb8c3igyimb61uaYs+yZWBZQdxBkBMzVR6V5JSvwqtP4hvR4AOBV3GJoTMKw1lenC5yEEQYuqqrp
jMqOsO47XHa/IecGuP7sDvvK9i5l5sZU8mqDEP2KnerpNSJgrTI7a8nqBhqjtkVfjx4jYTZuQGiG
ztu1oCBQHSLOLXOvog6Jia2tVTCO3s0LmGRmhH+IIPI3GmzkJLWZbjn/wh9qXcPTHGOB5y5KRFHe
sd1ae9vQhiu3ZT/z5NClD4S3pqIDcaocE0wUb3Xbpt/Uw+s6OkOUdgxdo57flkAzzkLbWsD3CQ5u
3B5F3xPPYN8ai0LB75JVPg2luJxF8t+cbRCoPshtULf0SI2ZEV8MU0ETF4lq5qwbooGmhPgNr/XG
WtNR7WMW5w7Yi32nBE8mz5wo6xTaMHLDJlsMsw5Sl8xVnlLHYwsNzc0Go7VVseJ3WrsAjSwnm1Sn
MMtyW7wj3rCtVp60INvSOi00Cw5yx72TSDDoMacvIfU3fpM2SvXdt2CoFXhuA0lhdnf0sgfSXlyU
PenQ22Zmr0T4D0SDX/Hn65OCGScBT0soN9LSwYO9LMSXqA5Rcz41H0QYfskG4+vRZkKMeIrYr18U
Bijf6myc7JtZOoidw4Ik47n5+Ni1dVruYgXML0Nht6L01aDl+P8XsXH8s6E+fziSbgmENlcfGivD
8Pw/Gjtt0gjdADjJ+43i0mYad9VTDHEsREC5OUTLJKITt+8kQSChp6kJvmncnEzbEayaSAVpr/Ow
BxWQi6rWMf2RfE0/Cpme+HVSNTa+yGK/ldezdW4rwCQqwSb/DHiqptDqggRhpipfvxHz4NID183e
SYi4nAD6wZyv1r612mPzvpPDhJ/aFH6V1/hUJ45F/yaBmRlofkMu5A6ecKeH/mdDVrwZ4cuXdmfy
tRa1A5ZgdgFdcWO2+qnGAx44tYhq9/DulTTxFba1gX7juIlJXshjWxJm60m5RB8SFZY3Bypq38wN
S8weDZaqgk7f+YqiBufjV9RjgsCBXlmynDHR9drZx9/Y3aATVVY2L3i/ffdInTQHDebsJeldtRxb
bfd1amUtc2bsNQfBdKahbpzguK6x1NM1AwqqmKJ6nT9BOxWL/KV+wGoIXXeFGw2H7eRUknSy3A4r
H9q0ww+NYf5ixct0EmjkLXK6+Vpepk0gp6OK6tyxS0DADRbC9/EVFpkREJmugmm+jKrTpnMEzEI3
+5EPo0SRtAwGiQ8s0ShDCXK3iaLGSqrVy/RJ4mm/NwhjsV9XrxHRsi+/CpE1CqKE8JI+cHvdZ6M1
d2P8VV25TfIPJ/A6wAE6Qu+h5gE0qcD5cRpT2BYEYud7gMNIrgvyeTIsj6KVMrNyrOSKeUtWDJHp
4bA9CV/9gTAFQFHs/TEL4iJZv66CjMWcOa3Awq+6K3BvWbv7kMVXCx45VxiitZwQw1YghU7zN8vh
wfzbk3OVy6APnleKNaq20dKi5iDGAjYCfXXRaV6z9KDEkwGslb6HEJ8Ix0Bl4b1X3HAg8HAEDVgR
h+O3yvGiUjiZJZW0cnkBfQcvGfwQBRbN/f8SDnheI9oIPDzehctmQuayWqwTAU+1D3p6tNaoMEJE
1PIxxFHWkOBmlwwOTEEZMksfAb+rm1Ra7LjWGcBAD78RCMftuFPlfJlUCCGtJhOPv5cSpPNadvUa
nEz0GXrejQhCB0HSYWXAjlkCtEKZKSUDKTJVp/Xlrl9JQCtq0E+pnIfgtRFQs5cdDNylG3BQ1Nws
YipLcM8OWkWZY8yawsMxphBsMstwMO5nmGoKbAkDWbsQIzFpzafRA/TVztDBEIwrkvQCwIa6pPMM
rkG23+fxCF5cYsH788I2vN1BacWwtQdC1Aofn1upTWvBmul96f4d2WaDuFYWfU5ATN4oohXT5X5g
NXup7JphOehiV8m6yKf6z5f8gDk+6q/D/++AyGCB8QBZlqnPIkMem51NEMNnqFF32aAPw19KKybn
UE+myuMCANhDrHvHeZKq789ma73UHMXdBThAKrHVs9/Kg2u5jDmyY5EnjvFyoiK50A0SvLToCTPm
tnK41BpyUjmtAMsDbD4p//zqN8Y5lH6tdvfJQ9BPhbLwBB8f52dAZOGmvd8RA1704tqt97jW8+0X
+NaYkTxlABDyZkgo00+mf2NB9NxtdDZ1kMFwYyHB3FQhgUg5Lvz+4syVgzVHTdWrHBiv5TpaXX6w
NDTXU6KhASp5SO1tN29ek4DHxsJschu4UFJrkjzA7/v+jWM/Hqwf8nzbANTEjcRt2q2oKN3Iah5Q
7sLJxj6tm2jQcU95I34epZVUVRwO9DFkweafe7xWyzQ3ata9nu5mP16h6TrRWVstN9cDCa+qIA1B
APT7qJL4aLTtKmNj6D+reshFzXFAaocswRO67E8tP259A4PdQAKdpuT3LpXFbjacbvS66EVhhhMj
asIMwpHRxKF1SiNaRAA8DxdyVWurJ+aT6WQfKaot+U5Wq4KYd1hdd4vj2oTIuMfVJmv2iJVsmvPZ
OIj73kYh+Xt+ijROibhC7c8a8LpQ/ZWrDwqUkv8Ao7XHdOe8eTt487mREyoWssA2t9FpvFKBJQub
JT/DNrEN95lpdIwt5WmkaYlmuOgz6dJyb6TO3UwtJW0yC3CIKFSAlz7Gbghugoz+mMNzf2CAhJzf
bpj+SQpRdO6zbEWgEBUSpsMIC3HmLDQOAMk1SVBkz42KCzSUbcK2ZfKXRLJ7oeD9UuvTKFckJcDl
1WiMZra4nF3gX1mU2Eqv4V9kooPFCMI64wprUIC9Bp9ZcrV0tkBR9WWGmU70ZGeRWCwvqG+knuAY
qR1eoZ4XjYl7yRfhrcQNutvFc8na/4kCoEB5+rLBd6v1X/yETHS7yqYZjSZXDk9AUFKob6pubPcQ
IdB4UVKXUCXLKrja1R4XoQJjBNb4TZYr+dBJ5++uZGGKz3QU+YziCAaF0S/sHyIteuUuKGERae3X
HnVM6wK9N1VRXqEX6GPcxp86Y9plMK65YojKhhEYDwvPg9SGmA5ix8PB5ax/NtUVlROWme+ysTZq
F9c7TT1ZEwXyPbB8IcZiI9hPmju1VBKmBkIVhQirkJlM4mRIXVV/3e6ZApkbTpcqAIU7V+1dtDwI
+V32c9/TbG0SToLsocGzhiwM1hZMP22EkPT8AvZAveLgPNsNkmhIYCbU2j7U2j6BJhl/UiO1YFzC
8iTxywor0e9WknunHLdbB8vO2bWijLUQNausOaRARYoZh8jX5iLIZJhCOMV5F+TgEukO+4yKRBgh
Q1q542GAs+0SP458oWmau9JrvAfL2jhF6zunkc6Dj91S5gz5m5XUdnRhI0ybdcS44lCHxGTcwmXj
oVSX7TdWoalH7xc4bjqs7C7MqYedcNiIvAADLLcB58rrUqbw/9ea9CBplHawm5Ao+LaUVbeswXVI
Bq5yMTdt5F54S5Eu2TDOM2fjIXmBdZ+MfyxBnv0bR1SS1txUvjXDgZahyefvlJlQgErBUdcZVMd8
U84K2lw9zq4THfuB5PGDAWsGGc5iIQQYZ6tzOSWP1lKpcUoPJzHC/JtVv9kmdmulkLgWNRSfRGBm
C4IQZxkxz8AvcicuA6PLLas94qs+b3OjgDeoQz/iHvZjG4II+n2Mk+nqqY+LVxJ8xwhlvbzRnuYj
SVmLUUP/ooYy/GslBPO/B8+FCUW9MrEyC4Uw15sdT1QeDVdHy/ZkdKg1gXgZJiMkx8Uc8RSqufPw
qhGg/tz71rwKGwRpwcN3u+aGIqI/8bRNxX7BY3O6Uun7oYfzVP/D2mlcixxF/ZYrBxlexXUXsJ47
XGMJqGv+7J/NEtJFqYmMm3eJRloMeahcXmmKDh8j+Zals3o7qFQeJxM/Q7g8wCFV4lSulEreV3r+
NjDl0axjWH06fNW31zTB82mG6vjz5XO4mkwCg5I52QHclN2Ao35rEoUpxGSHtkh4JxXsnomWkiE5
sJvekAJRUyx9WnQ6GywB+ND5iMiozp+BOvWYmG0uX1Cjz2aZ+H2UJRVFA1ZIl2+6Z6vZTFqDaCbT
FKCVRh2W2ui7evs06YejdldOGMtOXj63UQx0qXDE7cjvWq+T9M4v8vU/+DIRfry2qheRA9tu29OQ
aK4PXY17uS4ELQnMRvWvQpT8hLRQ6yo6P9OOAMf+P13JS/uxNqL3knr+06hL4hXhi18UrvGH+TyM
A1e/BQhf+ZC5/0gOUKpWLtsIFoAYRY711GpXeTrr7ZTv2g6rgyjPdBRbarhQ0NoqFjs5nfrW0C5T
gof/51+L71CrkbB+l1dyoPFCwPUJYc3fa628XGJwBbuxMHPlgRX6k4CDRNXj+xmdxjdzD9UVl1iJ
XVnoVheTDOi9h9OKjkdgWyQ+TumVe4Ca7y8hokHiSF61DG8XdN+AAOqTPKEmWT/Z1alJTxFysJaw
oSEL3ypsvboANST05mCocgClho6GJPk3vQXLlrhBDx95EqK72PEYv5vTWsF/+vZnXqNQ7Kw+TOxA
2NOYRLObnkIrmAczzrkh8lyukeTfuLt/F1kdyU1INxI/Un44KxkJ7uJs3JjqytrJb5J1HCzX9kyP
Se7TQdxz6GmbawzdrlBvqVoAIcumCJP5dhjw8JOZdCWSKOIZkZliYk32ajre4TIlqM+iO9YuJ6yU
aiVuAxl7oWo95EPwrwAOlSCn9kd1xWDywV85svcrwaXU5mkUNFEfvITpOClMpS8X3/X+3xPfOPLN
DQZ5rSfMYGbl5TiE9VIWxSuXrWvHXBJfFnMIWJSU3z8rhfdH/Jt2uOrrgbA1Fz41smLmNM95PyAC
KMtqAR21fpDksP4VDUY9EBYGw+8LgRBEREF5GQ31UARr+K+R3qGQcVufdvOWHAI3vTgdsi3DNO7E
tEp6gLNxc7ps/etTO9aR8rQfra7ZuL1+HxIXrHNUMCk3l7rYLaY6a98qnLnMLP3P/3yp5N82CgWR
LoMKshhieRHvHZED0KrRRkInWsHNySQeGPAp32vlzCKNd42fA9QsITlYlvG2gvEl6LpFouuz+1Hn
lqe7JN1s0kprAPLqLv1EYTqIJn6nKCVOdVPa1e0rQG+8y6kqQT/afupPi6zkgFS5yWDVpKz4El86
WU5Tu+S2wjPEum0EIaTIxja8794xQOPxZxmZmnysRgHAcN+QNDNwHqcMHVJfdf6HANgIOFdvA4G1
u6o6zfxMAYp4iIrcsDVVVjnUMfeTnli5ncrYWA8L7ErSh2kb2VXb37JIQJLaI+OK1jbnzHZY9m5t
CAV5AyoDsYWrkRTAncwMex+FmA56UwwzbERqiuISK/G/+ml+h67VzrnBKupWjPcy9GOjBFdsbRPV
pU4dO+VUm+x4h0caHkpI+DNNVo6DGFHNp0WR6/jG475MZKPRL6x81zeOeF0r5mTs8LVjyaLH/GBy
CLiOYUz2p3DPXjZkIjdgHY/vXNsnCWXimEybNePm4me4Ce9dKCznbQReSHS/rYUJfd6dysrGvA60
6U0uJEXr2R9K6flve7eVLPHByWc0O73DF1E2gHokdQrgSKEXIkZ1AnkfGk17D4Lkx4ocrwTyxoBF
YK2Oid4t1iJNyQu0yjT3FweCCqo0E2xE1WMFmI3JDpK0o6Xxj4cwcxf9szRh65zWpmRbcXGBvWXc
Y02btgcmx2WMhhI+Q4zyN2Ht3d6+FU+ALu6Mmn8m+/uOIfqWstav3izDnBg/L5z6wbV9vEEx7c6z
KdvdMMkhc3L5btTszNrsgsSQNCpu5YtfxoRezxRPnr5QhY+O35mlv6/U5OflmTaH0qrW4lzYIwpj
RHqyM0w1EK9k2Zu2F7aFK94EF100taon9nkryABphSdftMtzKdMWD0IA7acaVtlGGQz10IKvwagz
Ox2pZSN8s+g3TWofcfAZMTTU9x0GYV+qaTYLQ8qs7St2PewjSW/4n78mNLS5u4hC5QuSmCS5tFsk
BP3lOR2yFkF4bEbBD0pL5NCe4DeC6+IBqA9s6Ohfb8k0wgyTbSthIRFPNH46PsqOhyt2oi8VSSu4
+w3Cej+JD7NcZgr8sn0DGhEXbZlIdR5itxMvisG7vJGYizKEOS88d43HrBN9YRUAMDINKLr6wile
VC4AljKU2VDkk2fZK0xQdyOWUic+3VrZBdGRhIz/rx+0Rj9vCrM5CteOKXcUjzT8xu/hEfwizcCv
3betglQjvI/LBZA9LfXAaY8gzZ2E6QceuvDBOPf90jK0qL4HL3CFfwPnD1EZsVOxGGjBygKRRhP2
HDY2DDctlwGQynvj0ucFQKWc/WmhnhrAPtctxPzjPLY2qRIFSrdff6n90xSAOnESx514ZbHuopoJ
3JUkVlhuLxMpC9y2rJjIiavTIb8KJG57kJuY48Wy2GMmTDYpR/2oMJ1M+mFfZ/1iYjUQBNi00fvR
d3LtR28MXj1pL6o+Za7UeHP1t+vEwJ6xpEmaUjxxrcnjFT/JtWismwwZVet9MWyCSMLyn3xSAudS
TvF9iMOon4Acy9zez4ysibjViG5B5SqMLT3UlculRIjh2Oz+wnuyioDgIVcU8aw757rvPDwySabN
tnGofwnxbjfEvWs9YLRvdXto0yQv3jWFvZsOExqPVqJl/roZFjENBHaEAqaOJ9u6rbCipjSweN2+
MwYZOv5QHC29F8NToUsgwpW4nhMm63XEMncAPUnzwW6oQt3t75g/fGUmyTFOVkk9wAUloMpcTd+D
LGGs4UfKoEecve5k5AIHbeTAzuMmnrrZ9xpH/+t1LDxCCxR0TLfsmzeNvN1jzQZpd72rGueXhuBB
j7bqkZaoAEgLvSOHyicotArDqJ14PZHHtZxHxMBcdor+MDmwNHeeuVauxjxzW5KRPSKzDUfK4xWX
B+C5fLxqGVbZAY1YTnlAEDuyjBYbu6fLcaysVKvySE8Lan6izQiD4nEVe7NHAXZ4o1h37bOTvolb
vXcasgJzWRm+VkkTEwsygMy21qaG5EyPAeVtktIPj3mHFOmc8+aJKU4UnanEG053KfIpjQo1p3WT
enraQ6rkVhKXmYG185/X1t+SPsxc50+s27H78e/pvGT8YP6m/3+2tL3WeTdryvsJyV0frsM2EuwC
OrthKoWDE+KW3WKi2nZlcwEu9EJhOLLQ9jQ8sXzMKOj+JswXzTai0dVbZlBT/NmDCKHvOflqkxQt
wlBN6t7QBv2GrawjN+9JPGWT87PAuCASkl8QQwXVGpL3Zn9Cwbbu1ZWfvnBTc9PW30UdtIn8OwT5
FYy7Gxd+v9/qIv44NsePmNDRLRL2iRi+PWRByVpvAFJyEsCabHr4tFfEh65A1auqQVIiER4N9sIJ
AUMeZsMCU0NlZ+EIcE7vfS2lJQD8ila3T+LTsTA0OcTWKd+iJPU7gTkflCgaIhYqT116KIckLe+V
1eU1qhk9v1k/jS2SAree+Zn21UgoireNhkSrKmRm6SpmAjSCGR3Xh3UVeSlZAurmbDQR1hR5n4uN
SxI51vEZJNI6yPEbzHjKSM1U08Jz8iROakNgm1UkmDEpztsH5dU3BDOcCmlmNUgCUW806jZeGljz
7DvnuriT1G4u6YAmo96KFtiw4Gro4QR4gOaqCUodr1m9sQ/ruMMzEAavjbZdbtzUCEcCNjYYKpw3
XQgUByTCpiXgNobdLOm/Grwml19xeNP2kTaGCC4HHvuu+tC9g2h8IOG1Xf8TEFt74xuRae8h6SVJ
Qx6EUQx2+9SgcRKZAecALqQF1a2ExHzbx0uhQSqn+YQ2XhizxpG55B/50mUwNliy3dldSduw4eb1
eRDG2+5LLOj6mPRTmGg/TfGW8o4QQiM34H5wWU8ou4tBLt3yDv5tfiF9QZUbdh44wTOWlYEe/Meb
YVIf0fVMJV0OCDVpx2R7ui98yUPOm1XTjuKPJ8+s+PXyWFmUvzvsv26aj2MGxYxlJhHJi24TrVxn
TDxSZOuUQUjcuVXH45ACnkxYV7Q2ygKeNVlzGnVFXQ3PStwhuRrY2uUptTqWJV00iO8hxvrO0Uz8
yXxlHbmKTiYUDapK/VFcHmtmEBMGmEGz0FBV2Ib6WILh7l070vwgwgaURormg8Bkeo1yoOBobXal
5EBu8pQFjjSTc4MxBY6tnPWMf9H9xjDFobEXw/ZbP8NCNTRX5vDnDrQkvtd88I4mJtFPB5wOVCoU
2nubb6xUmusGMDBKvhT/t9UraGDj1sOW238MCaHA+VB8naYT69XPjVjyoHbJmbpwftbBjs1c9U+K
j6MuBdLqUB8heV0ryK4++OI4J6Ixak5+7qEcD167vuEvUjQw1n9Qo4uUrd2u8tuEDJiMvVHmCGEQ
UFHoopL3L1GPB84gXih04cDxlem5pf3X1JfsfR47rlh+BMK2xDKLqghM+bMKbvBFdo8+RQtNykdp
Oj4OxPmy8Xs1iBFDD/E2p2YqOBpsEfhRdDxqpWEvsfJ7WVMX9NcswzhC00cUJGfEYh5de1f0XVaC
FpcFn5I+hdb+p2nNZ11rdl1Y1p41Vc9ip5hQ5vVwFmWJ+lb9MJtuE/nPS7YRJE0bNpn3Soq/R+fa
i2KXSbC5vrbMvYqxv7jjYu4zxkir12A2B0TG31tCKXuvqv32XGT0kjKKwlxp7YO2t5Qg7/9r9rHy
ax+2Kk/kvVdvhfQd09NQAExprM7TgSfTkuJlCaBsL8jFSDsdQKg6lsCHjrfpFBfhgAOaJkJrSuNd
unrvKlBqPtgV9MZAnCcR+TvxOlYB64YFwqmXlyyoZgYpYYUZJ1SrZ453zGrrS4iNiZuvO3BnTRs6
KgwqlSTbcOSXdvILBGn/IOTHyMrugfYtQ99mSVBIDIdpMPtm3b8NXbi2k5DsysDdqzACTIwCqkSd
6kqW1aMudkYRu9436byD5BjMCdoIYX7neFe0m7J4RXfRaneiAfSNkg8dxSDUPickFhstAaU6DXdZ
y678ZTUS1W6oDOc+Cns9afH4bm25/0WZBAzJkC91HkTLXo5fJOSLQL9DE1yNga37Gz8de6k6zmpf
zP1UEh3kWWRjaB9gnqjXebBo7F8d1XY4HBHGsQecXUrMCaAOwYvrYOLsyksqoQYuxdrPw+zjjV6q
es6hLqhalDZ5GFRGLzROpVHCaBNIwAwNiTZ1wR8WKPJi2XWaQLkeyjWbXmgUkcas6yp6Qxy3M6DA
BBE/2e08GYr+ewsiPnmv7FeXIDCwIF3d4pEtMW25wmRKiKDJaRFxawpqUAjzuoHAGkCA+Z6wqpBS
I/UMs4ETEVJBV7MmQLqm8ARIxG8RYFZ08jQOrkFAw7JFOSllsWwsb+Him3DckFxLigwnxC68xKN5
gsJKvSdYUQrlozxiez0cP03FnARCzVr6F2CqMNlvR7PF2xsgP86+hanu5lz0LAGscPZC9plLRH6Z
M3G5cVgWF+KlDAPI9TpusvazFHA74egpNL0HeaPQUj4wJyZdV3ccaWJRug5/TI/JLEGF08joamCn
JoHIMbd7BjQqjZnuMj4PfUABaFvC1/JXlOayUVmVyRBknKT2Efz54h7xH1McR90+gSyQBEBfpSt+
XMz5IoBJT4Yg6ZumodTeWl3vVFwIkFPrxOAHrwZnpW29EPw5kdl54xPMPKO/uisiQWU+H0mA0zcQ
yqUYr2e6un5a3bF9frhJa2pPGOmHzSRmeu0cTX4XzblbK0IgYq1YZxRbnH7KMdYVUqhIY+ZuxZPq
UYqf+KA2G0perFTbt/SKtHaF6IGV3IIMusa8Ot2y82qH6XfQygoAOzkO2EDUWSCq/5PNbwSDnNb4
8yYB2aRtGesbAHdPxU08CdK6Ui9MwvEXJhbBQuhi0AkuLT2uR/X6Ln+e08qVkA22f5MEbtPU5DZh
KX0cnlpRT4c+yCPrJbx4ZUSq0IEh4KfjmH2DJC00eFeVqhsZrhsbCoUGSGxq2LC611qdsZQ3+suc
cFRtZfd+De2wGeri4k7ou68t0w2ZDWcv2aQhjUFukyuKuJUR63iGfYMZ1rm4KW2H7InYeWSSsxGy
jnbccGY+mbQi8J5euVL7qF5lcgG50cqf5Pah/5vdKqotxAoNc9m6qmj9exWpJcYyCP5G6Q6wKAOc
j379pMdGnREHHVY+6KI/Ztvqj96uJUM/viHXqNmON8Rxh64e4F7TwFnY9Z5WdhNDIccv3Un/AHml
5mrIQ5ZV0Y6i/U+AoqWBCclTUMzn//bzG1mb13SV5xWnS3AwThjdnpKaalF72ftAsSoF5csaPS6C
UabhXAvbmjNEFDqQlLePQsnIwLR259ef7KLDXDvGxBddKNM7/Nd/sQ9L8XU0LJaHVz8GAOSmVVYM
aqCrtF4whrcjDx6ZvHgEANKqakQF8RuOfaxjFg6AEecRp02u+ui3d3ztxNBr3zBRIrcKNm4oppSn
xRznvwc/rlwORL4ZFcO+sb5ToI56Awe0pUn+e93kaEUu15sYy0PJSXRRoUVWxd0DBpRletpPEkS4
mRy4Qrv+7V5XDihisGfz99VEtnJF1jDTHkjo2rFARNuf7rfEcyulPfl9Hq/3fr2VsZwi7xJ5MnQQ
CY+ja0U1gtbTfGCAKLvey1r2C5nRAYoDs4X3cexo6pO48BMz51o2/H6iSy98V1lHrmEgpCGbULuT
Piv8OifpL/h9LR2a3fDY8ay/xVT7LBOWKkY+oD/RkMM5x3m9V2Sc+wI9lxgpNeJgjSdWP/pAYCPK
OmWtf1osFGiuwaRPOdRxQ44nMKpjNMNeV0BgO82rDnOC+XF1BYQ73P54p4jKXpvTwBKwSGweWOXU
rlbjp4dMiQJ1o4Yzo6zHHKdAbTnVd/yEqblIYSL+nf+6aJhTegrqGmhCsFxdiq6TVdkDxfR/vKHs
/RBJNKRjQzWXt9GLgtH1pXyYSAzgIk6zwOxZxd66USdemTUNGM9W7EgSXf9ATSKIvSAtv0OwKEQr
kxx9mlK0NPl8+WfV6bS9kxEv47gNnkI2+VTvPa0hIv4f4dsRA/gx4Byj1faoUgsOKpLOAIibg3LJ
oNwYsxKL5I/O9boxzFJWoWo8u4oUSs/XOG2KCsgG6CoDAO6iXeBAqBHf6xDwFIvaBwOgSYaVQtSy
fyTRYxOrN3UtifEf4CwsMNqQZk6adc4d//fGimHX09NAGAtE5ZmF1bztpxbor/qUHnVGuhZPQHZQ
LOoJ9pp2M/TUzqgIPdwB4u5sgdJt5ZHC6H5HbhYM7JQgLoUntLzsjKnLLZMYj2/4+5WITaqs+kkR
RztQcbiJb0JHZmxDtpTOmFpdcUsc1m2s2Skj4zisKrbEFQZsdttvgBsl0JExrz2WyhvMjIRVZZQs
ZfHKbCT3tdz7j62rQf53Mc1UPOg2jRqOVBIUkcOyOygotCUk/UYcvX9I6xabkcJhoyTsG7lcateU
XFYG1EljlFUTFBPYZKJdZWeoiwCsXCOVD5NBNldPbni4bSzqaIYwJtI3wSXPhDKFibJ3YDT6puJj
wgAPzwu6TXMNC97iRdjQixva+zoyLPuhp4eZbuuKfadna3u7XC2MSDucaeOpd/nN9ZCCCnMxQvc5
yxpqvdU2VQ7sBt06LATmWt4rtBUp3kUnkz+ryEnCuUSrFTUgZbtC22i0K2jCzms0Eh7HCrzfpoTA
zyo1TQCatHk6YSAXlU/mSa4wJGDs+QDAg+pSONymqdHN7rEDWq4hUAQSpEsLpe3cS01HWZgc+dCr
c7qsFdmDW7VKNCSdWAKMEiAeUsbXp27CLko/NDbMVKbKN7xd13wC3OLxTkso/X9ZTOBhcq0ApWYW
wgpd5oRq3s3GiJiN2VYxtWlaIspOFkOkjp5Q8iMX87Qm+md23UvLUJ4DdH5W46c9WHuQsvCAdovc
Buogyqske3cBsNuTn7e7UHEPeLxZcKHqxvRf/UH9TVk6cYWyRVeR7IzPa+QnBby4ViV8UOBjyk/a
pCCEzCjk+EcaBl6UNxr2L8ntokjgQoTrTnKKIq+SZHWSHEARQxypbH6pDwZbUR8aR4ZB3yQaAmjx
XV0fA1uZ7E5kRADQMYkdxnDyoUnQuNpvqBBFNAf9tFfkUGU9rtzEV1Ga68Zl/E13VV9h20B0nM7U
vecmjR+kWllR322D9Ed1KR45XsztOvjxGENFEfCtOXpYEniQLrFpba1GfyyRvgKK77fyX+FfBzZG
UNV1c75KPWjiefmLc70azcdOnNjGxFYqdlE4OyiR1hetyu9wEaXfdoqx7wtnDOpSeelDMtUk++xU
cxcGVDcvz6+w1eH1i5l68Jvnph6OHO9slLibFqHShR3XoTDzW3oHaSri4ntrDjSVC41VlmvwNnSZ
hzzzBVbCrvZkPVyNLesafILUO6Z+eePwQ6pCB8QGtQpC9NP7IFKvmy1/5ZjqVzdnn5MKrzbQz6jL
0q0BjQZb8idvINPWe4zgVYI0FOgz6CKRpf0PBQuLzA5c+ZcpHgvbjh9JGY/8qzXwl/PFCdr8mIru
JhpdMopRg42hPDIQ9S9nNyayxFCONUtMti9oZQ2Y1grXEyEkCI5eN3B/Gg8v+krQ1oVNvjEC16F1
nicAMtHSceV83ofpqGPUuBLi0B2cB9szuTjhP6DfT30wGehHr80jbjmjRPwRgg9sCmidaMPbFP5V
SyTRMLhFTOEOgJ2hGWZkpTqaBfNlB7X9h2paffpXBeC1Nj52JRyJD2Vkpq4y2uXwvakm6FVB6FqE
gifVnd7EW2/kvpFYSD4rguREbiEcz2MZJ2JGp7KDb83GsATJzRh5Tx9Y8FbmEUGH+s4BBQ+YUvTa
KEurBfipd7XNK1Em7xmR8ErYyu7frua2PflheZZk/w4VW9EyjqUxy1AmC2znrZWvF5PG4QZr5xsE
LLWSkVd/fsIgCWjswsGdBbU/C/J9cZAV+1CCCOFlBujcaRVCWAXUWcUV2HoiC02+VTbnrYCk+vBy
XmOVjubp99qj5FOHW425+wzGv40e6krTzOEEvLgMpE6k8j80BNoBkWtk0xULiw80ib24KQEMRw3y
I2ZRywkK/Cvn1xNGTxvHCgzI6nyaG9U6M/dCCEBUVsahnnI01nB0ujoY0jE3RVO2xXxyadSM1S6D
bFe/EFWAJYkILOtmQVZogxRYGy4V345ibJhrsjPhtL/NKwnBAD9VllrxOr+r+oyCsB6dnItHNvji
N2FUV+P+o5APvD9SuPJnghfElNpg+GJ8gZYDXUXutEbqhhRn8E7TfE1a0vT+7LGeIP/rIKnmlzly
tz+JHZ5JhuqPVR5YsawTLlE3FXRsul/TpzmHaMmlocSb86tipOBdYEmqik1/6wa7TRNIXDcKFpDl
ZA2aroC0Ij+TwwPEYtqyTZztrFavvjPv94SCczFLeI3L8SltFP50xHQpsBfRpBzL7kW3NmwbLzWI
+rp6c/O2J1uF6F0HK0XZK0tpQI4kKT1CcUkaCH1DSiV/EeWS5E2dsM/zG01OoImyd/UMP0oEA6Ys
2eMxuZ7vR3C8yZlX2/unfCuYtcOLfUGTR7NqtQrPmBDh3+/UJqaB5yiXjqYLe7qa7OAFy+H2Oi51
tc5plKwQc0N/wYpk0ZjiUfaK0ouzVptx7EXlxSYrvbtK54DWJE6Nxh8IoOo3YvXuWmqDaIS09iJ4
7FUDm6Jbjsegf7xBbS9W5KpsuQglvHTfAZWJtLsNzizKLbulv+LoP/GALrmhe3r3R1hpxZidAM6V
U9rY52xJO4vzt7m0CeXM67+Z/RDnsy44/AkQVWT8RfP/3rETxKjFsI3I+OcmjRc5YhJSfmZd7Q4/
TKmE7fCpKUK6XjaIkwc5w5vsG29+7Rz3S21w8B1xL2/1Jd7AIrUIA51EGuGgchdbo8TVTK2s2uIH
lUoE+Fa1HDS/P53Caam2BqFapN4gkCdY6cAglxS3f60Hbj6s9lSMZBUvPiUhrjuaw9uu6ivLQj3h
cZ+TlD19aqDcbqrTiUbSNt+KiBhlvrEI7dRI2rfd9MK+Wk1A5QNpNtg95ZgvKgAuE6kv/vq7Q+iY
VgEOe6YvGW4g2TBeRqjS4F+3ZSsnc/VFDUetNlD3jD5ItZM/OFWmRNFwiF8uz3wzC0xr6r6diSRG
I8s5ejDVcHwZYFvAjf4u/7b8gqDnQjkoHr3QJZx4GiUGbTpvaYhUx+ZoS0P7k1arhhVlqYr6DBeX
Ew+NN7TVsRqCzUEZaCtQou1VB6rMLnaXTOoYTfEVb9Z9IJdeQKYaLB8x2dqU8YN0j7+PBoJycpDr
Hy8qLe1qLt7ZZL7+ha+Wesdt7ytJoebqB/LMFViveOCGCG3AK9SIDNuiGEXEd0O/xnxgNkzNkJy2
uB/9wlO6kVtnOTHPPh/hX3T/AfekeQ2a3zciGcGFuAepC9bzY5c7AXLj5w7omVbzNsodlqGUYXb+
xwk/YcGa2sUjOwEOvAVGE5mxGZKUSqEwxz7/n3+LSuqfnkofAVrmYKx2a78rliqXcXfZp7hIr7dA
EvOLSYoasONE0ZvY2yv6LaQgnLZOKhoLCYLiuk0sotxXu4DTRBigtcweVUtkze5kWkhl/Nz05BQT
IxqubGS6y2S2JXNOYCkzWRL76HLSNe9pTJet4wl7D9F+TnqB9zPc8rr0Ln9OpFAaeb1PA+Vfcdqv
myKVlvugZGVgQFHPzEZWunayM5YMtVvfxRumPJOWTOdgms80FMto6PRunzp54y6fcH0Codkf0hNQ
oI2gxXS8sBl+24lfH4TgRZpCLlJ3XHNFUPpMVvNcwKyFS883PIucpR1QxQ9F2Rd01/Tji4J+Q+vC
5MfrSWxjoxuKBhcXG3s+F6dsji5S3P3js/FAj6J/SlQsVvWs62VH4IPSJsrXj/FRZZZniWZGF8s4
UQW3sZoLuB0X9nVD6y30f6CdvLPVOpQSMY5X30yPSQd1XBnpQO/mFbae0/rN57MU14iHvpjiBTr0
SqqHyYgdV4Dl0NKFFgcYELsvc6d3YALnQwxsq5nT8G0EYhJr2JRn5ZKsset3eVBqBGgHgGJVmxNT
PFNAg1+d2WKSW0CSwp/zZNH+BL2Uv807YeqaLm2CA1NbhIkwELMQHr1BH+IVnWewHTFO+HJSMYzj
EuI4GyGG4Z/nlu1zKiwbDxdjTz4NcvxbS+V4qWJpq1OpJqGiy/hZjxOj4RrqN/f0wtNZuqN1DoKU
HrDw20lAEhwcjDkHw1PZOJRVcuSgCqhTXaPTEnCBPcP8u3byBts9y6DFU7ffIRx68lB8SEuiu9O3
xOTg2gSnICBlFz89UqATjWe7SmnIe/lZnRhFrRhb4kgQKI4Fzdnux1m+m0I3/sB0BbgLZUuJKXhO
M3Z3X/we9gyiWb7FXl4akN+QNtw23M6VfvTkaRqVNBme9lG1sdsla3d10vK3ij0M4Jj5LSiuhPrr
0FTU/x/8+x5NldMsgxuX4l0Johyl7FeTlaScYy01R6rvEBKebXXhPPgOWf8KpmG4cUfOx9NE9eBQ
wuCtQTnn09xUZavamO1dqK5e5xM0r9SP333jYEaarlO4rh+AIlxyVcvoIovvrVGMwslJq4CY9+u2
kCYJCZuD3TGo5vGpStPxyzYN5w46WaCGkV/IN8gecnEpB4N2eIInCPDl5YdWGrXm3K8w310GsKgu
IX/rvZi3yQW8yxxK5Ci5SptFKLAEyNUws2iZo94UgxdW4TiQitUYgCpB6SlbFLJMuzGY6r03htqA
M5QLhK9FomrdTaqMMMpLazIQ9Ht4yTKQwIGa2m2A2iU3T8fhJJqmPvb23JkdVvCCLdRz2kbBDnyr
3Cw3Z3triILyyTV12xLBoo/16ZHxE4PXuWicghg60S9udXbyA9GS8UiMwitLJuHJIkuU8nocQ6fj
9UOQcF8tNE+CaAVHBP/sN+biCrVZ4srwjcfdwiBb4Y8Kku4g+nnuKTw74tnvWhe8zQYwGlEPtTSP
wydZydyfOMWAAeF4RwpK/yvxlI1z2qt3dU5zn1fy66U3AZSonY+udFQQgZT4mJPypVIkCtc2uvcH
NAZpLL2wUs3XbjgZ+HVbaE6VfPPgzFvUS3UFdIRPzh2+3PHvpXGllCzSxJhLZyqNUdVd3M/4v5s5
tvBPhqqmn4mWYastJ01yTgzhnzRDXFKFwqai6w/twobKeEUswHSjv5DG9D5ULiOn7NL1LjLamYkj
tX4IA8jif/t3QPb/5hCPniwUc1M2ndxjW56dPEQNNO0wDBum5Kc4QOr4UsoLTSCzLLsOXwyhA5Bw
yX+QOvGJvDfifWk+K1woNh8czgafYpJ/Kt43VtEj0UikQn0xwUYvDlkcCt/SbvSMHVqTMcOP77wi
1hZ2q08Y1MOZW7+Fyr9LxlwlPH+Oz1nmbuNWPWOW1sEyWuzV9fy4jyaYPS1TGoS5/oFFP+73rbXO
dWn+4Fv+/kjL8B+T7XPgUqoGHwk4I/dSpaLSP61SRLzoRmY01j/FWKxefElZqWoEGIeh81MLTT2M
zHXj87L4kEIYR2PsHH1tY6ARHdxoRKAjIymj1XkmDveG2Ru0tGaaen7yR6ODNgPP9sEe7gtytDnp
pAH2Mt0k5DfcZVYxXKW0Fvbb0TD7UxIEZOOkSVqnAFr7ztRkwQUHQ1vhugi90m6zRLs6iEoTXrOe
tgA6MJVLeeoJcpWDlW0B0DSZ3YGNKg6Z32t8YJl0Qc0FLCuK+EoOgo3TL2QjyNobBZKx0Rgb0ypq
egUSWrEQETw6AtmxvqigBPLeAXvoNawYbpDMtyh8RFqyjrtzKKhFFPvZRQqSDADs1UQaCXOOT54x
FwPYIbheDOlRdFgzMjQ1kJuHnWWM5riuv+qzKEkA3jAzKFUUAq8W2hvPUa96AoS5yfkw0Lj5C0Ey
B45UEsGltY6ktgawETP6D9ezDLRYxKg/C7UO0fqrxNE187FAH41mryz6nISmvcpFpMrPRUlkexrV
01Htpackr0Le5TTvBwbGICvpvzchFLN6hcA17g//zkO2aBQGq3/2tseta5Vya7NDXxstc2UHYUtL
EX2jvLbR9NaeytHclB8FmnsWArlMFOFR24iU5Dzk1iv5ahMCs35GphGyLaSqDbDpJxrKgbCZ1Xvh
wD6hnqjCJKSEHNE7UarTZpZAXwUtnKVz+Hl+nRXvt7JpTmSriIHxxKTB16XlJK9Is6jKTEI6fEvl
fSfK27O8bFQUlAc5jDLa9WA3EKgLCmBEF1T6IQplvx/r87zRh+vHek9KjNcX635OMBnyQ30SYK5F
yi51BznlBp4ZbGWoPNc88NUlkvbkmI1gQgtvcGSXzPdPVPLo5bkrhuT5+OS9Erpki08HQMkjxyFh
URa8edDpFoNZYteGRGi7I6sv93vYslkuwstK4DpVQddLztMuIZgc+WGyAvTRtVGQLyK9hKZGeOWP
stzXvIKrkRRsQAXCnAWwaULwFN2lZXRLwP7tBe3z5f16IZY3UrYaWV9DrSgCF/+0zalQ1TlFAyn6
UzupDGnc7q9jwBNgJltjAxdMTgqJkVS3v0YVd4Cp8+Tu6Z5gpW5/WZc8ohqWbk2Hq6QyMI6VB1pX
xj/pwH8RcVcD3tnaxQIH4efQTh91PnQeSE7AYCs/bQjCXONccPgwMp9Rg+7Sz4V4DEW9E6SUr4BM
dhVF2tEJPjc6cBKEJAv+2OGMwNiOknfxLpM0ChH2H5JLjJGQSRCt0nc1er0k0np55t/PtBFkThYj
UvAPVAM0X5MBFbz6kba5o0/P2Tg7Ygn/mHDXTE6OEggC/qB3Y/SaC8yZEXD0z16ZeXZo1vaD/Tc0
YsJky+dmnDzIH+oTJU7aY6yX1XL+y/5GxSKUZ/CMSKRSc0OLDYq/3m6NFd1jVIW2J8d+BHBMaR+N
xxa790iwohcv51cj13lGI264DMOviOFTsK6AlFm8GBFh1dnoyVpqpfIhXC1RMROnez8+lKu6p0kS
G899pIjulJnPsZrVCOqbvUAsiLD7e1nWCX3NIF9ik5/crHzSsT2eSG0UZy9rBt9/611iR1gNpUFQ
5mtTVyX85gq/XyC2FXZt/LSBbAMetBGAIjbpM1MqGla5pf70plj2rFf9bYlJI/O/qpIldXtXghjS
OrDsCA0U0eK8wmdnpvEw3vTwLCshGR+a0lMGi1F4vX+n4jGszUODWXyhF4o1BQHBUva0RcQj4cs7
FWlRZMOt6hOZWH7ucRzKFy73gTUyrLIlDU2/NnVzf2tvo6l76OOSr/TjHuoJOhA6XhqZMoOiMhxe
RVySfwd0RxYX2X6p/+6PpYoatJq2G1scj4o3CBlR8EheZ4p3ArioxMr4WPvg/IX/wl18oI4Kn9rI
69wjbueJ3qK1QlpcNdp47W8Zf3DUaFTPXosJYj/LoIJBrsjijCtuks9EP8rUiyV+4jRvCBUo7nts
e8K59fnEAm5XQZbK6KU47ECh1lC7+SK5ATu5WluovhrdRvOdyKHui1DYZ87dk+TZo+wtQaACjDpz
Hi9ckba5rgLu4nrFOiwX/OFEWRCEqstUpALSl3/Gd3krCRAEDWQL1aoc8CwjPtP6zj0vbon2Nmfe
CejSgAQeYuOKLxU81d1I1y6Tgp/ZVck3WvKSIreQNRHLmhd54zAYmFJ2XOBuIoKmZI2mVJKEEcmV
NiVbvH5jvp6Zjjzozvzc/4kR2HpiM8mQXx1pVqrr8UMRAEH3oCpXBlQ4HE+xbcZqj1eMlwQVWxZo
8b+wg6qT74I84uGgCmayeNLumdLP9aROFcTKhm03VcCGOFDgPb4JD7vTZxlmrwh+zMqc++0f+5NA
RLGq7RMiGFLvktI8ohpIgzmJY6IZeqFhImRdDpv2s6NjmUNRx0v4OSTF5WLGaldjblwskwY/X28/
8PBYnCCTI/DjOSmObNc9uK6bkks6pcPZ44zvYeCNU/fbY9DwtVI9YGYb6lePabwMWEnApw0Xpf7n
vyamE/eYj1C/GUIMh4e+QVow5hH7Es3QApWTTbZlvp6fRooTVObpQgSHfPxBLM1toXOXEm3auKRB
X4D4nKTUgftH74k7Jym968jJbctCjFPlsNjyEscsVLP3brRL2XW3j06ZBnIS4mmQI8cwb4bXBhpC
ARDsKSKxO5712mW3izNdVCh0ZQV+8uwlorwuWeUHG/G0iunAPQhlq8cAPW3t2iIeDMndEGdWCg6s
B1jM0L2D6XIqMqMwzvDmYnuQgUmpV8sy4TRwK8M2MECbVGfpcxuTPeeob5KYnA6xTVegvzHt2xAe
tmgG0GTeUTn1UjcwjfYEHkN4GTWH9WCT3fsGcPzblNen4SNwMbR0LmewzkecBXRZVH0FPRPCnyx8
LxaeApibCrq5Flz60JMtpf6SczDM6yThRnYeFDx9FD3TVGuHQkxA1tzHadf95b0zzOi/ygPGf44Q
+5H+N6Iigmkx9IeAeJS/i5zT8aird//vujzGFUcnps+P8mHZFDVT5pR4HAwGpaYpb+d8Z2ebJb+S
ljoR7TX7EwkVFtMcwqLowDjMFeHlrkaMS3TFrWVyT8h6tChRFBOdU4WUzm2278UJgpp7s5stq1q2
oq3I+zPDpXAerqdEyqW1D9jCaNXJnnY96XoX0PIB9nI/cPJqqoA356mFKL+ZG0WMHU+anJ7wB8t2
N7X8U8FPTo5jXmMJrPRS+vht1wcRKm39s/Ymg+6eQCKtOe6kPBStZ73+WRfXMrrkuMjKRFCvvhRV
JnV2xrUgIj5b+qU+pC0a6x9ztz4AIlHF8pxFjOa35wfrBZ4qPu2EXPmjdg1wAdWUZcOuEUhbObqD
EKkpUsdOY2eclBpkyE5Bcn0a2TQuLruFKR5Oa1hOTil43g2uS2MQSuMQmdtTq2pXT6yZTQARCk7K
l5VF8GAkeAk6VbvBuOlLEDC2ZCUhM6fEt4+VmCWIHgYYdgfwjECA4dPMk/FWI+xthAyU9W6h+TFO
mOXD/gqsSveXH12FhNGwBuCq1CO1QJheKCmi0OF57TQnFrFcSY8/JqqN4FqiMAbEdxuiPTwuAEwD
v+1S5o3ZSQGb5Xkk8jmgY2zsIW0MtUMA5fg/e+33NId9jYNiM5PsdzodOIKEh/IQPpAMgqIpo+Lg
lQCQxFa5i8zSQ/t8cOGt+mvbtLuWLyi4cDD1uB0P1GKLY3EWkOP/4txmVngI8bt+sRN44Hpr0sl5
UeUhNY3MtZHRkd7xMQp3LtoavmY+YYDAmq7cyYv2GB4CBkGVV7fTUy4yffT5jU6AL0QAejIOAQKy
4Yue5xDyBWVIBeMNmoCUvSfc/6qawqQoXtxp0pkXdGa/XWWJSvcSP4NuYInee8HwTmb01/g+T1Hh
I0GxsMU5FV0cPIzKbcbJz5/AmwOhvy0lrFodt7dvzxfqyGfXwG0zsqXlxRQ2xLAX2bFyX1skBy5o
1FhmV/+IEgDdN+/PwztlAqsThSFFCzXDQuZp9WRuJKWrUewQnYo62gf1Q58gYW+h3OJy50GJ1TpY
Nt0fbLcjjBvUYVmb4dCwIjCpXUfqyqK0fUSFsxcqygQlO0N4gbTdHX6d9rW84TFYF2PULc2NOetF
M8IGDuLCSYmgDR3CEki8ax4/4RiPuGQeln2BIMvVZtAJqKY2LKF8Zq3gK1pq4FPHq9RdWEqL4zt9
5qSzK++gqq3oAQ4YA6Z03dItswWj8jDmtaEIS78GettXN+yjb7C/WGP93cnbmsZb2909enGZ7G48
MOtf1/3kcExbMqMCFuuRgDy+24slCc0f11t2um3M9jnz6pj79QQvMmruHeGGWqBhRXdj+bC6xfh0
x3liGk02CtYPkkfcsBLcaSxNLRKO2cPVGN4jAJNUQu3zvdFe2tOtHPsPqF2JAMbBN15S5fXzisf8
m5rUzVODyyVSdNJvyGxGF10XPw/LaIKcXka+ICIF6qMPYbRTguNnV0E9l2Ag+kEA+E0WnhirPrZq
Kah9uoZDM/7mckMZLR6cnOK6uXVSzbuUwm9HqgnFGM7b0YSQvJyOCB2pirH0qIZDg3/1wqAKb2Ig
kI4ZhVl/vlqnPEDT2BQ7oOc9lCQ5uq8DR80fO0a1jn/hhFm2qsRE46vqqzzrbNkbDqJpduUaGsLP
6wf4Xb+tDHc0qpqw42RcaFwJnHgNtQDJCK04pxA9+dVNQyiTcX/65iepFgpHCxWtDv47/GJG8jeX
YZSDHiG3KZ5sFHMD5btcjwmFbVjgGrTqf3u9J9bZqzSCI5wZo5cBiK64bnopPUlOZU+C3vuw16dp
GOVnIO0W0oQ3pqBRLZeZSIDKgO+mj9dwNm7TCFp7GyhBOZ/ThCUQvaw0L+soNKH2tafwgTxUDW9k
RY846aokJws7WL8ijVAXA6hXOqsnLTQjwCQgHi3JW7ki9D38W6qjBlKEbDyDSUJxsK4G75BPiPhT
BjZgGJ9Z1IA0SC5SGIlUznkVpXBRLjNGYOBC/Q/wkbUK5sdfIez8rEASIxOWd5gOIskv91GMRPy0
rMEq6BzrnBaSllYXZMFEF4Crv3MGorvWs+Z68Qlheoz336nzCP+anI+z/9DfkSjYpnew+fvHfTjW
XbRePueZIKrJMV95wE0MoLhqbzp8qBzESuF7splLKGoAKoQ7jN/BpZaymN/0+/EwGGl6Ut8yfyHH
3GgPd8Teff0qS3G1xOqRevQjUeqIFQjEMlPza2h8sjmbAXZRDr/1aasFWmKRy4wbk5iUjnGpTHim
3aZUzB+wwBL2irrCl0alNz2Y1+DJe27a8hdfRhB2XLoQ+HZny9C0zw/rvIzUB6xh0aQ/1uX/umF7
BJd6gfYGsvQalWFe43D4QTEHT5Lk1d3wKo0EpdemvHBiGqm2Fa3BQmVzJKpuWBxcuaeBcalOG5sq
pcuXHU3thWUqpC9PB4hv8Wx550WjF3EHWzLTzgt4NFEx/Zhx+ssyiGHf4VVNtCGG8p1SZMbvMp+Y
Crzezohf/jZrhfal63SEzT959zTJ2j2vFGOm0PtxfJfG2cIOZcaOBLoH59eF90YYPJs84IdLu35r
6HbwK95rE3//gC5t82Xn7hIMSl8zJsR2yCyY+jTajre2ynQiUH42Isu9uDX4rCVPlS9TYu/bOMeL
Mu9uympVovrL06iNVx4rOj0/vtXwQ2wVgI32FrdiP8bBMeIFMwDpsKWqgvD5H3JCAsnvDYc43k93
eF0eaTsYbgfRdSQ3+r1hRDM3qf93Aklcu0496WD/oz3cU1H5UYQQOb525JDbCIUmVJfnuv4zUCnd
0DazModzJNutgqPrvpnOXxG+OgZIbHAPLkyn+mct8faqnr9b6El8omrEnwvdI1YgXlspVnzjpjvJ
Y7HBiqW9biInoXu7bArwuG7AlZMJ1cptFUSLtL6MXfzFjpMc1rGT04jPNJTOBzJk79IqX7o6czpy
WXp+UQmW1ZSYD+2goUUaKFostiZXJdQSFNb/f3cSxPDnAGii+ghzB5ItrQ6VoeiDQbuFpA2azvbR
8uIzRisBcZkiHkMXRU1z+r+4Hy7KOlz5gE1HOBMO3Z36xYHzpHhynKr9Vhq4ZHz0U3HWKqpn0cZq
QI0hdKu3BOEF2xjdJRKLNbQzJeFLNqFmynnPfLj9gLODsA57e30kbMQsCsi/DKnhiqt/FR7sqF61
F8RSBBSEuZTkkMrG0CKE01YXlFRqoAR/8OgLwCRIj7UZande02lq7P8Az5fXNF5cVPf6Vs/NnWs4
M6qZtjXpgyX8dPKcN7d8kvXxSBS6EyiBCO3yhSLD9DvGOAmVffyxgO5VO29pbUllazDTiAU69Mok
84Vd/zxbkJOesXGseDAOX3wSyK0VxaizldQGxO21IHMmzKBRSZeIuRlBFl+5E8d2/vCtb38KSRsm
F/ptbIWuXHUgwrdrhnXrChMQ/E1IqGTAuAoywpVlyYUazRclT8+rte6aunhyHVzRDUXf0+oFkJkl
xk+yMRYxscjiXPIqVIv8i66L+Z6sjPEs2OOCMlLT/8u3hm8uvuNX9M3aOJAFZe6rBE5XVrTp8jbl
f+qlsDIJVCdmiIMiXQrpwdBU7GDrEQUFyva+jgezkrz7MesuxrIqt7VYMhM9BZQpWPKyGTpq8B5H
cURICUZTVriQfN8OxJGnVUQg+g5LI/wYHHUgBWzYlU+u1lxcfVhG3J9e0ZbcX8U7+8UnZl+bkdKz
i3ql/52ZyhzXDQfaq/rwk+apW5k9eRKP32ZwIQsgYPFdCQLN964HRV+qLm+4FbAzRtaLjHV4xmea
pEp0shAsFDk2E1HX5zKsfNZB1Lq/SinBeK4Y5Ql1dz+RhkouxglN47k2cA7wXfWgz7hRUnhbPfjf
NDP6VmMla+V7NyeQ/R664Ul8PMLNFfxByKE39smCLj0eg22LSzHaoLSDETrkuujAVTQanCji3N1z
XE3czip213VT/BoDyuhtI5cZdxc37YVvo7kKIiAptfqnZygLav84YUfWnfde6cn6w7SKqvPKLqHK
27BgGfMgW9h0E3N7jKmiQs01s/XgfcXq2T2Remd/2DTDH0rOD9SWEX9iojj4yUtyFTvwpuQtrWdk
Gj1VDRYyHEKNrNOrSn7drcjGmlsxjzBlLzAzuHDZVXUlRVOgyY7wWDl/1bNMMEjfopzKYnHuW1ku
N0jPFJaBW0pQcfUlnwKNAx/VBp2S4Ol6/rE101qqb121rnsurVH8V4o76l+mPDWI4bclbUCBvGa4
qO4l8bqxmEaJl8ohy213lUVHVcXzkqt7tLVrelRs8NjhMMrs7fNaOKO2IPNDSbwqSEXRsGYwhPx3
vumhA2wkw0N0gEUAEtglfirGRBuJbLdG9DBFmlqhCBxUJsBzlQNh4H7HMIX93buSY4NIYS3iWo9w
2L0CTczDyuydNj7Uz3UdEn5KmFln7vE2OVliLjfBOGMAQMvyXTLQP0StSUmotffAik/aik2BxIwG
+97ALRoV4KYsuzT6zKPFzZmgS5x+FqLCdG6lxsiSI5+vyuWJTBc4C3cRD4slVsd3VPavR1F7Qsi9
brwujve+bAS/F2BaztaCHliitRO6MwTpHtVA+AD34N/LEtDAMPRaS1g+kdelvIcImfMue+i5lifT
uiV9zghEDf+COg8wj0LQ9EgF2axYrpF+spcmTegAGcQJd3cJPkiofChhJa51Vtr4dG2M9S+eqZDv
WRPS/kpAlCK5pTy7ZBgdvpiz0Pckqx/tMkPSHKZ6MGNok1djQRda9lpIxVo51yr+Wowc9URt5R6v
6TiPAIpqLdVN3Kousr9VIghlBycjEnS1gb9FXjbTwELcCeg1MEDcAyR/3TuE4cT2aMdWjs0bYLop
G7rauZ3QHDoyfK9G7kHYIWvosg+SO+4M+WSVWVnn0GtTClxR3grsmbTdQ8QFqCTY+aPIzLmdiYUK
nOgskYfC307Ka9gQijzlQ1HER45/EtDRVcR1mj9OoFGyprKD1jloFN8mNxLP8XAOdqcjz57xNT11
/fpuDQgIbrEKO0YmXOuEKxVuybX0LYag3rJzmfRNfoCw0igTo91TDj2pFGiWAS9uhI4B2GjfYuLA
c01FTEh39beOraJGE4D4eJQ2Z1HfvgsDEKH4r3fXknNpR1TVF7PSFJSacQmykfMTZdY5NoaNjZoJ
FQl86hePXT005JxAH3NkS6z68YCqu0iQTKvtRzavZROFXcKIiv74OKI+RwWk4cTlftrz5vN3GG+x
EO4+4kJSnEMWGaFirjQiaxzNtf8gPfBz9Nl3DimTroil2ioXrAG2KNQeP5TMs4yG2VGL/roE78Lp
WlsjlOmFBx83xZ2t8EufdwDY5iSNUKZcsU1/fwGQDxWpanj2R+XPrj9X80PBjLHiGwrLkwIQC24R
xkFUz6RXZRHQr2mSGhRW2A638fG/4VO8MrTMMfBDHRITjbceW7Qm6Sw1Xhm1Y9y15KV7X42mQ8Jw
loCQ5OSGEeVeKI4OBz5wusYnq2MKOhQVGTDiPy74sEsvR5WnnoweImiSlP3MMqJW62mcY2mtGx5b
XKc/rRZGtFUKKJFfxjNUe1dg/hRJc60OJGMoJIvE/LanFtA1bo80tLt691Ktb2NO97xwT2eTrwqk
Jg+Hyp6Xz6wXTjitNLegJLIyqmRf3JGIldsDiW4XIL3EnUqt4HIAltx/Ztmt085e74E7TqiiM/AR
Qm9YHXr4yGibLkrlC8uKRwBeFAawJEUrkKgu6wN6viZS+6eb98eFmqJdyPJshL96xeGx2z9K5Fj6
xhNBo4RiMwVcK9FyzUjxuJBdJWZtxfijSQJelcKwwRWxmoJJ/Nb38VnQELj/psl8zPF/P4L/OF9y
eHZlVIJvLgxKdkLJPKjG1gQl83bedpmTrlEqS2ukSRem2MAyMBi9coIjQn14xrOCbAekKR9Ibucb
Myk968El9E2Uo/GqBpTKvPHGZt2NJKXsU8DSPbx0BVAp+6cdZMMzlMUsEXsIebKODewhR410NUmA
UBskug4BPyseKB8335FvtpJAodTtsS34ztHmAj6JnB+t4zMMC/0C5j8029FU+ZqUCn0AU0opqNQH
dpkXIg5vo+JpBzMwuOI7dG/oTn/xceu1QvETis0vTRqGnh9sISgmCHIfx01DDOKYwfv5y5E2SVMU
wsubw0kwXisGry/Br2gZEKJjzRSmS+H5v53OvaV5DAfWeaf6Ou/rd+TcyejzAoWnkOod/9lhO3m+
CEjtWEkhHlhK4tuItT/L7Fg68YGECWpPFE3sI4U1U7o+lrINVTcUItMFrim13nlgN5ApwK+Szh5G
UXverTSE1MwjCTMHuspbBzFjcaq2TTxREqYfA+rjHqT9QXWrTpnjF5l82UK6r/RiSweZDBbwq7qu
h3ONltDf7tv4LgUcg8sPEn9y4AR5U1Lu65Hpq713GMIaM5Gw6vpjBkDtANqzWQwQ38mTbKy0QdjX
MuWcCm0NUTrXHeW1L3vv5mgSp1rd8qeGVg77ASOCqfuYWKFoHbz2JuBY00cHSHr3p8s1sKUtfBeT
tiXMoLKMwjLi5bqN4BaB6jA2ezo8/oQfifewIXNl8rzP2dKhtTbgQYkWdNmRTEi40s7SKPOJfZ+R
3PHvKDAdRpxCVxlTsdtoP9Eg65PWXsI1yIZnDhCDQvzjzU7AbFu6jZp5Lh4x112iFVQJwCi+xBgy
EAozztR+1KDgFY9FKo9z9fx1qvn2262gnKtHvCpod6VFnx44wOA/zG6c+7hjuWMuz90S5F5ThZO4
jYeXGLf/B3h4CH87aKNOQ1iFTDgU9M47B09KjrKB2go9wI8t74dG++KkqSqGrLMazpELQjQHOWSH
BnEXgZ7Afen0HjPPeLXdb2cIhW2SHPq8+PQlXsuFJxh3bypDM5vDygt6XdhKu2E7ZOGmLw9q7pOo
DphPWghWW/9OXPAdADomgz0IdTtiCLCYTHYOT1qLp8/91H0RM+07tQMWr9RXZe48aA3EZ0JG36ua
8PmwuU2Vr/b7XP/MW2OaN89k8DOGGDAGGgpoBPVESI5xBzC6WE3Dx5yG+zTOf0BEblsYJpwJRHri
tHG84eLarKteUvvxnwP8/8ISRoMMsGQ/S0KQ+0aRApQGggridl6ldO/FGqUFwdDW60xZpHR8YF6X
L+e8E+WlM+7dMiTAdw9LQL1RDP66LCr3M7DdChol/xK0bFmStxNPeeic1lWfN5sooIBW+BFowanM
IDMqSlnmRavfuSWfjqeE6Rm0sINGEBTfIRcjSz6JcG0spsQQiuiLi1nkJwl2GXHB/ZcdDLw+tq7q
A8Jz0cGcfX2s9dtKVdbqaU3KYLyoTM3zliSqirlsut2VyDsYrHllJ4pBWzzpvRxKeS1wGR+ahO6O
jP3qwOMlYhf047d4mBIhau9MrzkC+ekl4wNn0IGXssFRJqFYO4Yg6S/SDlkGDrCHFgGnSUtEDnGc
+h95dia0UaeitaYwv09mfe+k3D0vCjd8C8WJXMUrYlac+/c2XaZL8ZRFfzFvdSWw3rLE2dGkNoA0
6WzgGvst0hyltlW24d1BvwGcllZl5pMbRD2HYtvlVJGMYHxoXM1NbOnPmXdwEg508uRmuRgXp07y
L4VcbqXoRNX+bx50gBV3aa9VgBixSCqp7B4kCJX9mOMZMmj20T/Tl7Z4/3ffBXBwu9Tg95JRph01
/7pKnMltdI/LX1s9FsTKNe5miaXUI88h1jWiN4TJvQ5Bwv+68FW/0xYqPm5+eYqH8yAH5d3YzzQo
jBsX8LVWBY/6AD7GVxdWcfabKN+GdFK67BYJcUNLpJLy88B/Aod9j5rhtbZ+P0lgccYnk0AHpc9R
chJ6GQwTpbInHOPkxKR3Qq6SADil+jcX1VOWC5QoHeQZ28bR5uFCrt2clJS9APfpRbkG9Zlba+HK
EaSwcPR4irVjVM0dsvT+7UmH18zXRKBYJ9KWce2EU5ctHTC/AqdxDP2QeUivCy9XSTHkKRJNjj6D
XrRI9+W0hTOHak4OQccmhYW76EQpaotHZZNPyfEwSPOoRWJt0tKl0Ila3gueXQqMbrc2vCzbv8kF
ZFp7TL0VI8eHiary8hKscreNlPWvfM++Jj8QuGZN44RAR6l0slqyyVNMTULitbuMARbliq1nzpH8
tPYADM+GdwsOBA9wqZVQMDmia1BfCPq5Qfk4ZDglVE2s1byGnlhe9ts0nVIQpfhB6BXat0/eLQ4v
GRj+Mzbgt2zNUXhfgL4hF83sjSnqMgjYyqhfIdaVvlxsS/rbdl126B5s3PPJLdLIDjXm5MhPR+1d
g/R4niHGou4PUBZeyTGOBof258LygIiiHw6U4IwdiQKuNHrAgoiDsEmASaRf82tezMMmp/VkQkcq
mbCLHouBJLo89m36MkVvDgYEYJTnCleqZ++EQAHwH17pXAa0X4bkHi3k8dvYCFD2bgRCQ5juvafZ
HZoJ4IZOfm8PI34OLhKN2FWbi7XmHBtOV7DN7pXvp3xGbD+ZlTUkLwRNFh7U8IMAlBql/qhdI3w2
re4DYVbTpmpTNGZDEm7ugm4Z0vcODYJ7f+dQnxNRtYU56V+L6a9PLbPNFHzLkMM+H5+Mb2Ew28p6
mM2LfAZrCSNgMuxuX/YFWh79G1htnBDr3cwGKY3TNv/Cvnvmem8RzUIdwX7Y1n2+R/A1vdeCdgxt
6WNMil/eLotn30QHpOBScdgVV8jQ0xMsGLgAHLrECshx8SM9+1byVd1mrwC9uOD8qxr6hZMYIB4Q
Ewa3xVC4qb5+W/EfUeiIO923LlhetH2hsyLNel/NuVCUkHX4JoC1y+LcJURgbKhsf7PepBzElxQS
EJaz9mjrWq5RYnIECFUSrNvchatKdQJcFMn7VwuF8u5mci+BeF7wBkFycdzUHiD+rmkS0d+ZCmhY
W9vMUfHoWrX7bYdwDfH9QZ6W+/8Mkqf6qp+YEA6/wFhW3NKym/6Opi1qxTNHG0RUYSSqtkMxPXe3
G1rO02yOmhZJD085GmgqbAAd8eofz6JbF85bBqwXSMUaT1+nbe4aMr864zn55giyASWt/LJEhDPt
o/vNyEnNYQrJiz4nizOWabYcPDYqTlYViH5rwmjEsIHfoBG66dkjUELId3Z+GZbnh/Lu0RLx01Md
8y7T3FAJZwWpNmb+QHyVdPWhZ1IoqcgIRszhwa/O0pU0MHb+BkyUpR9tP3Fpt451wJdwyLoA+D0D
objPa03G1nKqJnAftzCYLUYOR4FOYc/JoEHbSWv3NB4hE7ctDWt6T3YrA62dHx+n2M/Ob7l1Xcht
BfOJu7NbbZqp45J1plXk8JSMRxBs08nmDSZ5hEgeEobJEVl1Zxb1uYjZEcDTfvmdS3+TlIv153TV
ClIAJ4T8Ad+G9UVHnMpJBOJNxBbGRReDaTy5E2uDT3fDdxFEzxd+9QvHNwiEh4P47+IdqK0BmPUy
6VcIZa3rCV/xnfHJTbooDhygjQN9TnOSVYV5Ph3QVsqBdH6Z7HUsfLVP0OWQ6TknMNIpfsApAhUU
+YFnQN0uAqVSOA6CqR48I+N14fUfUVK08k6jTmDy580bynKIxYTUjmHgmaR+/4BtaqYITeoBp5KW
LyWZ5vXDnFdrStlISonXPY/xRKyLD64Q+EtQP9R4QXwOq7zHYOU8YrK4KFM9qf2NmnFtczqQ90fP
Nsq3G6xjLo2yBbEbhoSsX6S4f9EPVXz0pgGWbmdSdi8xT9bwU0mK/8VYXxnpXJXTecIH/PX7rnBa
h7XSQz1FkTZOgmxoU5q2XLKVuwAK7qhhCzpNTqqyKiKfeKtnwwz5O3voW1ICAEEvEu9jPHD+/1P0
5KNkMLK/yAu+Imw3j0uB/ADSoV9DTcUTf+tlaijJKUTq67YKZz9137wSZnfOJmYInh2H3TXT9CWm
nrXLDMjsJjbSrBjM7ubRRnq2DSAoUGeALVABa5Bqlv4ACClZgRj8BL5WJvPC8scbpVaC6R9kljmo
ApQsTS1NLsgFeGec/5nxaeU0W3gqmYLHY4FfZzNjNxvSAQjfH5sRVLRf5v6oEmzC11CP2Z7BClJn
vXGIQel9WXKxA1l3W0VwCQNqF0nyeVFh5H9TK1tiOGcMY3Lf6sVUlYON6f/cvB3iT56GISr44gY/
NzUz57tANmfxvYvohxPYrrrmx0+5QK/mi23d/EmoRP67LV01696wjiygAWbBvbItS8toBJktNuAu
/7bZ3T6YeOcbIwbssNGPvjJ3R3A98X04r3ShhlPRz0hdciZ64JDwfh9Dhef9UpiKKhqv/NysKvpf
Leoo0SX37mNHbhNQcjCTsPYZSlc+GH8vds6IVx4LSQUw0y6W4D+M5UKYk75F7IDR6uv5FBbKvhZ6
lyVygJV2yWr1vy3KPPG/m9SHkQQM+AZIQTkYcoJalfD+sRZXDp6vSIjJQD8eIrS9T/aEatFXpHAt
cxrs2S+do40k7VQHwzkSElPaoAgY75Koe2gc9YpXZ51C/69iRXOy2Vjt0lLIQmct8GcRVXAa6IE2
ANEDSZ39gH4/bLoCeJia3MhFH3Zp41lOSLScELUhfurfOxgK5Rnggbc7vyRbahyjFVliWW9J3/ac
bbtAhw13uncwK3L7Q7XcT62rc0Ly4AbvODfUZQlehZEyvCwbTwoSdcTKunZzN4H0cfvo0tAW5X5r
LlJZxZPqTNHd5Kqm/1GBpaHa57cMx8MEwT7ubUWZ943Dd29m2He/2VFhg5BlUsWGxrUbiWoDWHv3
ZdGL7GoJBVpwJNm/Fsp0AYvM3uDa3CDO4xb4g0//b3Qc2QJtQ4OhtdlRZPFaK7uCMlaoWseFVaPJ
urL/PHiDbJ/uFzGj/7khfB3PeHHy6W81z7E12yS6mVmMzM+hn3Tf9FgACrR+WuI5HITRI0RurOJw
ewdJBs8FbsBnEMkvDWGl1sb6Ujssp8nvuva9JEL11VYI0r+duscrB0MKHoxBsnZRBs/vK8xsrPGs
SOyeyN+umIV5ukxJ/1RtXjv2Cg4z3Vdh8vqhv3kFGyo8S7FNWm65LyRYom8zu/MjvakQeM/hQMo+
EIjhgm9NiedSr+Ld1cBrF33Woeo1NFCJq+JeRjmcUy9201VR2C/3z64IgLsL3JMlDs1+rDV6cOHw
usjZI0by/NKzKHn7AZm+wAGmCVX9343y0Jyl2FQBV6WbtNBobCQvhwq6bCtgnwR6OwoyRmsNQliP
xVpfqYXJYI0pjunpnrrDIIYCXTT8PgA38SIZsQzg3bOtX7eo8Vuecw+XAtVHsro1VwbyUXjVx/Iq
vyzsrEx3cUvW/vgAjyZiYQrhz1ksUJ+G9syKi9UF3jaY+mA0VjFT1MtFTpmcnQi0WF9j18Fj/K7S
S6MlXhJ1WWExmcXViiZocgFkx1BDgNPnuwtf2LviX74LFl8JffI/JmPi8DFIHHz5Hk/8nSaqOpOx
+N5IidwLuzalG8Z4k0PPt3im0xDLgMNq6B+ubUbwaO3Raund7V5YboDl69W47wMTMZfZTNB6D4Iq
jlnHBYyr1IFTUJXyf0lAMBncoudzmF437QDxYUBf06bbT1VINZmJsOzvY5LNj2KWSbgJJsY+QFIZ
2KTu60V+vH5IOw9Sku54XrpREKczOQvP0GcMXZ7RbhwtJDmtoy0W7ktZBvydAXWFRz6qCCXK4u8O
b6mSjBkR3s3T1PYP+QjwIPgz8USZfTt5NCBUb+LAQDwzuQFgS0fSZnSpg7C59MMjbIbgqPmauoEH
kDSfP9lVJ7d9sTUVhAQrrmN4BKq2OiGD7eCRUnPnmGf/mbqWYnNvNP2JKYiKNF9z8xOE5by41MEv
mv7HkyrHetixNZpHipPSA8nf1EnGnN8IOVj2uqM2OCkHn3sSn3jbcHILTdDJQLZjYEz+O5WmYFgl
Qvk86p9CU7AuwrXp0JJyxloTP7sbBCMhQiv5UrgSiMdIQtbvy4qgSIv82zAlrWa/79qjXU7R7Twm
WJHa3ZAGX1w7bMj/iL1MEENGbVuuGfsw3Foz8bgY2Lq1s8T2jsBdVDfWeec0B3nXiQjcHN6KH6K/
GtWgwKaDMm7XZitHGpIJSj6Z151epXXW7W0VhoqX+eZWXdNe5WEOUzQRP5H4tmUSrj7izM7VdPQX
CeYeoIUVRF6smiAF+lKllcQ7cfSHvnbIFzOwueHEiWLn0A32MsizP9Jen7tndUeGHqPCvj+ngNJU
7FAe02uFtWPFeTzqEV6ettbNGKySGJUS/Ji63IK8YRWjC4PdnTaozKtgNhvTrY0MdixsoyBsI+iJ
ZBtTK4fAF0aPv1aZQBylPvaJ1HUb6E5ceCv3X99IrjjAh9kjN4gS64ESytCjGYYDjaEAV61nire+
lU1+fOixcVNjqDFTxX4gQlrfACYcZAYphfCzymHVIWDO/nd00/jt8lNK03+KpxVjE0Exh0BPXMuJ
BprkY5y6NS6cO8TnXvdWzv5Lbl3ISHx8g2ZdxvKAD9G74wn/2/7h6fbrYMc8Zz6OCF6xrP9gh3DJ
J5VaLNVTsxdvT4URTLEyUekM3fOJe1TzTuXdQRagTlLAHXkQg68Sg8hyR/c8lCbhdOdm+3RTjOIg
t2Hzt4737lT9VOUm6RGh9mknGr4EoGorklrNDtZXklKFWdLrgspjddFR9gMJ/KJwoULxE8Yaqq8N
Qxqjh5oMCfJAU7UFN6d9VyouP8SI9pVvJcf3E754bEJ0bCjUwdLm/3ZCzMRPWlMFzmtOwZAh+CHr
D+ivJyuwl4oaqf/mC0gTwnSDodjob84L7TN67MPPvVLYXYED/JH3VCkxfhd7+UHT0OAn+2KUEhP5
+poF+uMLhKWjShmO/6+Fw3ivTvWWYSAXYrah662dmpGOH39Wp7oovlpIaDWfKvwslzVn2peuMQHT
x6pkxgYt29VA/QoUFJ4ckG/Nfww2ErUb0r3CVuMhUgOsWTKG7DDK9kr4rUH/iTY9mxcUEKw3E7BP
QFE1//yoQLqmttn8nNtWrFCWDAbm6Y5tM5J5rqYr4iPaWgcu3rfUXDTZBtSZ5xSsR51R2qotr1qR
+z6wmG1oeR22VahHRY9oriJdj4SRiVBWXEdhBZ73Zdy3d0CIZNpFbQcwBNB181i/CJAsPZRWIFnz
y15TOVNiKj7rfVLVvwjWALWdvKBJkjCVRe1YmbBd+9J1W5YDdswECsFTCkNGLKiiw+PkaGxtk4vk
klVAkSDpu8eTELdyEhPlmlBCojQmoEcytaR5OHcj6sXrDxmoQ1hI1qtN57vQU3D0gPbChRZjIex4
JYCSz/OrPCjhzFbDn6ZWEKPLucWtDK1ltWQ6ExtxQHpzEzHPNP8MDBvG5atZcYImDNi614mi6GBp
q4L/CbMi+c7DNUf2PiQLMpZXAjPiNra3gNxVhguCiCOQtKIqTOzd8lq9ckaiiJNOXglTWMQ5xByb
Uiei5p8dzz27/DM0RAtoXR4IJ0BfFC8xJoKRJ3BD+sPBto/xNdyRshNRD2WhEcxAuTwN9SQy3J5N
T2CRgDG2zYFlJDuZelGKz0FDc9Tv5lxh8eIJ6X2g8szLhhpyPi9FVsvhBvmfYNi3VKHj0k6maA9a
MLYZSCIAfpK2GcLAHNxSgPE0YYm5e4P23eevnaFPcjlZuRjd06kXo1+TqF+VWq0VOaDIACwrPFCm
o1bWpz5YMO3w/vwk+OIAdp/KhBYpTxE6eTGZk+VJBltp+yr7bJCv6t4cl5zoM7k7uSy1CRzmoQW7
zjg+4dgMyKOcY7V1r/svC73OAE2+our90qujw3nGoHAGWhwCBvWBhKFfgVa+kbCzk+YavMV3gAFD
T4VsXAua1jEZ0jxv4LOAU6ExuALHG2oCAVOaeLgH9rj1ljgdgCa53Zif2nsGaX+U3DsT4imbHOmt
TBaoykauoG87xcS3sZ3kSGemN1PfllsuY4gwjBij0WESLiNX8Js5saH38K3/hqZQqeMYJAMD6sms
QGbFpGQjfcTf1np/xE9ZYLQQmTyQRSgIrgi8S6XY5cIOjtW8OTKFpPqdDFzNoOAVpw4vu8/baLIO
QnQqqfS/EcHXKwrr7YzwFqXiSHxJg/GvFJPNKhO3lk8Yi+yY23mVgpijnwoeKoVWPLT8jq9Kc4WA
+oAWDkvucbcpKfVkpo0qn+qSnZx+cDDqPW3e98hGeRvNcdbQgPzQiFhCj7AlKMZ3bxQqhiHb63bB
t8juPKcDTdFfX1JWOPiAjXemzctv8kuyE6wwtGIlWcaI0OXhMnXp9oYCOcf5YSqwcVkEn0plKWM6
HcmUcnQd9EvFysdJq4yul4DyqwJNrEEJG4S8tHx2TfHaqVzuJGRLuV+/KycMDIRSt6CoTCjlrpm7
ptkFoDKEn2FFHH3r/5VUx5jB7mz6mciRh2z7SRGD3WlSl4xqgl4yg3xo5d/uOAP5lai25ryR5hWy
JXCogbIHU1SHfBNrS/8aFWIe4MQLkwZI+Y8AboNDzdwbq70jFOwOPj0vKMynZ33MCerIG1JhizZ9
ZVbSiP0TtI64LCMYnPKiMbwIPomzIKYdKOIGATEdmQ69fEgEMAeICBJtDIFEPji0BCdcCt/tXbiX
zb2jwOIxfxhKG7klX1r69OIxH2dNWp81fT4ZC0AItQeG+RCAV2tbgz26TLEzupy4YS2WQTJehdC9
tOFJz3GhjuXbE0VR89NiG4O0sV+rlsckkmJA8KdDQ9mwQ5RYxy24hpARzHRePi1wsi4U2PghGAHm
k5bs7THRWastzujmHiEf9eeFI3sY+Sicgn/uVCZnSI0X9Vw7T63ShNruLhTHEc5DBytNcGBMyBcR
BKw5zDi3FaFUjRfBCzGfbDgx69BB+lHODWceLGqVzx6dFvU33eWotDkI3254Osr5cYtFeB4ATQ0A
+s9xsISqtjlLiDIfJzi6SKkNGaJXxXq03hIMquLLHPvYMN/g1kHsov9eclsJ+H+EmGHmMns32w93
roey4RIOJXGB9L8GvIlCO0KY0PteNbpnvhfnSWbc7VANbt9r+mXFRWdwD6ZpldhhNqyzdMS/sUSC
TkssWCd29/M+XnJMIVsRxMPAAWSKXqP0128oWkhrJIS0AoPjsWfLZkkYYv4SLon2M9f+YeDkVKw4
9wjZ8trLqqPnStltiO0S64qVAk0/u27Rf32w9ff2yRcW3iHOJtLBsx3WHcinhV1nYWBCbcYxGSWD
EhaInKGnSEQCRNeUp0qcHy7+Ni+cJTcqaRYniPSSYZOFYR5VuahUEoFjGrEnwXq6PF4whwYNTUn7
F0U+5HWlnc38LyX4LQp71TzUWU7vyZXN1/muOoaESHqu1Yyihm3kLq4kDrLxZRmTcmbbSXRxdMfS
JE8jAKx69u/QRUSW8nprwisVo96fBAchmDeUR6sc4Kl94Z/6VseAHeTs092l69ZbDX+/HCWCG+15
T1gjGhwpSH2bFOW7MJszBXIpNT0L68ouKB3qaYVlfeycBOFydsJXDazEYKNIC+dX6RRkPcy+ogX5
NwlT4K9ZNotx236GzmShOoO1ly/aAX+YZz/KFhvBH/HDCNlpB/gSQ1k1mlUkdn2wck9IMn70+0/8
9XRfyJJMCuH5n6WjKU6Iu+Nv7toHzr8vP7IFQwVLsavh6vo0bEjn/0dp2XB5EzvwaN2VXdK5H6o5
Hahy3TFNUcw/+kiQdNrbyeF/rAV4hD2dmvyLl6vV2Z8AeuAmupzzwcjPce/BB08C8fUzuGo++3R5
WrC+tdxaR4TrK5PduZnq6a/97LesadIX2+0DdhxylPVr47m4xwbjui4qW0pKUa/4eoakPdiigVyR
hGVBDO2DLjCpboOh7I8jcfkTAm/+j2CEfAvY9SjKFLbyvi+7GP2C2t2v5A7OYzP/GhAg8hSA9hvZ
1OemDomV8FIBgRlCtv+1KMYLBGKLeIey91HO1RQ2Pb4eSY34e7DXgGxo34eCibw0SE5IdkFXnbZ0
Fd6Hke0RTlsM3V3CGO3SA3vmfsH70rCU50wlH4HUa2N4CBazCzR+Ij/uLdT0ALlppCLKdgJFOHEn
ntX/QsVGFn3GMsgsBJFXlpCrO6tFD2Wjkhv95GgaJE3Y/vs0EvZ5/N/hE0diDF1rz5zT8wymax/f
Jwv5/v42gHI2HKf9JGFnVpgXPJYdfVBFppE8wL4QHGFJclP5Dmd5EuCgVAkM+iaBj+Y0H+qM3w12
qaivKfqjMJyU9ulJhjy8MceUB4Ed6lAWS0ugjRILuxXP3AiMLqNTmderq3GGM3REWbEUBk0jmRk5
1aI0DnJmCwYc1cI3HWrMYuej2LFbP8Np71psW8x1tRD6zOL5FUrkeSGgeB0K4dlGZTZ/okdq6GPG
MLyneBhnyJDA9M3mCQqlD88TQC2TG0gh7YtWRLA68qLGgyeLaLAxaENxUigxFT/2yFbbjbawrLpX
qHxU8leb7a7ORdj3WuOCCCh6eGWOxjZzE66IqzqhEZgIRhmsy1ve8M+I6ZqUeDlgfoaEEMeB+4T4
wfsTbXLTt/tJUjwYWKzGl+1lGaVdW1M8AYuAvLV6hxqh8AFRdNndNExIu0UNhreNFNkgLSaLcNFY
FWGhcvV6v3Jn+uSm6Wkf44BJKEd87787wmv4FGoTFxjD7GyV01mhd/yUbHIHYY2ER8fnKa4Gp7RQ
KphabzTt+eUER0QgkD7CN4+jPU7W+Ee98piaxztww3Lpn+YoTKt4Kh1MiOqdxZoF2UWzQ47tcBDC
VWOcSxZPfE9avRP6flfLO+XKCrb1u8VzB7qeoLZ86Xv/3A73c74T+ZbjkJPgQDmZxGzvXzQykbgv
oJA4V7dXXpTRIHQNU5F8zVV0g4KcVwldtyaKGOd7U9gXAvnsJMtq1yUK/fTXp0cL8aN/bk79V0Yx
DFYHN7ZuQ4n2Dvvh4s9/IJ55BllI4B6LEDu7qAtwajnLewnq5IZntNFq5BKmkT2heEGLSNom8ztk
P/F24Gz5W2rtMNDH+1vaqwXJDYYdcsmSzQ3oLrRfhL3guWEK7X+aGkuFPT/2FWnFEccdcQpSV7MZ
afCcFc4+qt8lbTbAnrhVcnN9tnxPD2w7Yn/+JMS77S1MlMGMpVyco1uJ7sfwoOo0Jx6nYM7L0eOh
YdIZP9FvZTfppIMPvJqB9mCePNF5PUN7bKUZIb9qG4GbSSEvOPaDHWOcmHaZcjqpKDwUiWJLP5mp
aGSDmw2/jNZjNvtBxGwjlXWVmAiZNeUjhEmAifhCEVOFdp0m3fkteCPVGSCqzkzh9+6tn/nn2DQb
7BF/Z3PT+1IsDxkn5dqGYTFuiVF/EDumgc+qVxXQ+qMvvB4hMTP3A8EVfKOvUshJc6aHQ+jOIUXV
dHaUujr99mD5RTnrmGM6LJ/TKmffMtodebPY/7aJpk13iYLQOn8rcAoeIyNV+HiMu3qkiCJj3OKn
OcjCVykt/RkV7V9azPaiMgHlTgH1zOZZm8xBPZPGyaCX0j+AZUn4EkJPk3ObLm6HgmrB6u/4SbE0
7eBHlREUm9DLWa3Eoe8I1BJEKbb0PulnNrKI2uM0CBYktzG2JzbhnmtDYAAharNFQSC8ZOUw3bwe
0L6FAPm5ynaW+r8cK3/v6x4kOTF2GS/npQioeKBEvdBZRGD2hraCQOkOi+CPpP/2gWJekUamYV1A
v887axs3bAHTA4HCjf4aoXTEVZ9I1G6s5NE/8TqACEad61bIFwY8OJqfb3YAZeeT11jsR6y+sawE
eNN+YRWS31rlaoZdKVILExkYdFc80dGx8F2NOlGQtlsJ3sHnrn/KE1I+FKemgrc2sw1Y84zV8uFe
WiAcaVGdTWPehFdLCHcRDj7VK83l0c0+i48U/utYZo7Pr1u4MuiJiDEh5pFVnPjzg5ogF/Thknbn
TfoACm8DnDSOmgrZpDbMh28/4+rdIhQuQ3rKj4BtqoX5HkMuuVAudZwHTKU8blwVeW2nxSWkMQ/h
yh2G1vhgD6RPVoPv6oz4a0fRHdR75pqIQT77UG55B6Er9K2s2wR7BP43VZcLi25+Uka0PriGfoSz
ByRzcvuiayiRzL/DQQMRnoUJQhOFI8xQdpDuc8cZBCPRiPT35/w10dEdk+SXgbH5AINho8l70+WB
GCPdb07nrwh/fMyqRBGiMDkrGtVa5dxQ+KxOh1D2L2+kWmnrTyronSB30HlklMyGmRmzODWR3LXm
eeS4/HCaYh60j8FF9nErTAh3y3THMlfwtBQfsXrKH/IPeLQHxa0VCT6XoR3zuUbyCddymF5hT3rk
Gzej/qTIfpwXbJFcoQMcnHCi2211QM0BOZGD257inH4JTDmJv0yQmSHmcyuDVo/F1zAMuaeWvuNA
1nCAjuJbsXhu7RNlAtKR2riSIodZY3zhNzPHCYuQi8EH7kQ9z4SwQfdK3NnoTg3eOaHoY9AMz4s0
ysBOv0Mbs6MVUgPOX0X+Tp4/a/ewDTkMlL2N13s0ijepfVVxc54dznK0BtqSERf1UV+ES+giu/HZ
Dt/h73D7Zy/U6TxHNFBCmuc8Oa8rZG3v2jMlyxJBPWw7ssl7rnRkkl9gaj5z3zCYFdc8MCYzBWZd
Q9APmrahZZUNbAVbcX60DcaWrCBrL03v9dnIWy9h0RNvZAyYl2SccuPIxR6yap4ktp0tPHVc1RXl
NGjhQX2UA6O0L1UZjcMI1Hi3jUXZvtnJx3QXyqT3PZG7YjVKZqWFaIR7tsIsI52SU8DF/Fnr4AI8
wA2MzTaZ0zJGMSc5lZLEa6eurT3yVvCD29n0gs2mb4T5UNrNEDz4YE3/Ur50LEJlfCyTbY/Z2IOl
tnh/Y6oqgJR96KMwqTfBOXylD4rixi2aiGY9ULr4YVbRP7q8GLAnnv6u0jWa4d96c6jmhAxj99Gz
Xta4MnG7PTYvEjch2m8ef9TjQnnv21MOS9lw1M1SwhaxZe1W8JCHQTY7ta+w6NzDA03FBr8JFovZ
TA6JybR3FEeSVdgtzMYSqGG27O2rLFZ/LrMUtbWHqUHDnnFr6ROPQaQ/Ph4uMvjLK+5IB76o8Cov
Lgn+0DKZPAsvs02V5/qzDa7oHwNJ3NA88kflJ5HP4SdMPkjsWdI5j25+hKGjpS5L6bwZLFcZP6Ab
PLWQlGQ+N5ByyzP+tUDuTLu488+4gZyH+KvKTOeph5IoQkSI66WybCcpKC9xIT5KV4aQztLkcVEa
kCLSKCaX8rwxWdM4IpTV4oFr+KnSqveRFL4nM2Oz3UCgncYQvQ3PJHcOc0QUUvg4RhRmp5k8u7bH
4Q5P66uDeo6CDM9AhCw4epGGvAoVmUUV5JGjen7heJ8O1fMvpSBPSXH2QcgAPDQDhQu9RMXl6fV6
A75+CCOGsXb4Of1DZHiagtd7apyqnRPVFG5N7U+WW1eBH1k1VAWHBf4KoK/UXGJhKvESM0k6cBsu
NFpExNI6bG3N5MYkZAH1tF+C5JZrat1TVLBervxxB7IB+Z0ROJzIa8ShYT3rHVsv40MEIrxbGNgQ
pBWAHrz4Gsk3Ccu07RutXPz4wvwsaqCV8qRzZwueBh6tNJO+zA1dfok35+Deintcv4XPDF+Hh6FT
7p7gRZQe5Ndid5FrYi9CDM4CZXkQp20p46OLgLKVRZfTRu8fc1hLSe4YVqr1s+1qw67bNiqeMt/f
bOMFqDsNGNjPL1R43j9HYdYEHjzPgmXxWicXzL6tgiini2iB9VQrstepboRt2Jyw2GE+D4uWF2ej
UHKZhQTeXOaVo4Un1qAR2oGScH2wci+VNionehYuO5yxjoPynNHHu6RX9wQUXAiLENNwrlhrV4X8
Y7eD/oVb9jfI5ag3Fo4eZscegghXGtSuxoc5qMUKFT+3CyXWpDEo4ZZ0u6Z0YkkE/I6S09XDfebw
A9UnN2k2yrHqrLPEzGDMDIPgs+2GSjNZOOUUh7hYvG4qbAZBL7dNG9Yl5eOujIORja/8useFrfas
HZ/U5KSdzSBTpW1qBbSATmX5tOdKs+fAC5Cs8r8xohkqwwGOCf2m3R8wrFF8rawWWX1yZgs7TEZn
S8gXV+AZCj2/5cfp60yXyAdTAfMmJUtesZTArlv+x+tuDsUYaK6n4K7/DijvOZ0IqURlBz05Pd9x
TAq4KAejW9nd3wIVYciUvrUVp5EVZw6h1w0fkqMvAru7sInjGCmpNCdpSEhEz+/3Bba8rb1OWZfU
gAOmBZP6iSohssw8SJ6O/5fZWYeSb27we1nM99xePua70K++tU/6dqEV5yetLcDAtOQg2HIJLxIc
FLnSIK2YgsmyXPfIZ5xcGfI0vZIvHDpfWZAAPAVpLKJkbcfj7CUqYlFaRKJvF9luwyB8GEtp8GbA
wSsr6SP8ayaHeRQ3+Q8Ij1SP3z8qubhsqY/CyyIiT2qoKkntaWNixGv1wjTIGUw2k/A4333Tti20
QtfGmx4QH5YiM0Uwcue/wTWRToidCv+KM6X9jDHHZOatcjh7sIq1Ql6giYwfpZeyRYRIn1zQODhK
xCbT5aG1pQQsufmOIY/RfiDkuiars6v34llpc6dd/LsKQBzbk9ZFe5T4TTlk4xcONM9QzRfA65z1
nD16NSohAafFAUUOSRCn366NugV/CThWDdD38VH4vL1G8qmCzoUEqhL+l69gVVIqL+l6KLchKrOR
sYRYwKCqqs1+oo30aN0e/oZXy5/Rl8g7IOdKDXvm26tc1nsx0DsJrQmvyK/9ZPDFV5mI4lgem5gv
t1ipGp/aFyjiRVRJ6FfJTG0uK/enACwGgs2U2xvWDul1rdNnEKFGdlyUAjnlxQaq1kaLS5I/4277
N0v9EYt7Z46gGkEOUHthC5YS3grRgi0zmUeZg8YI+xqj6iLpQOXNWK7ke0ulMDVBECbxUdIn+ZQ2
5+rA4JbIPoticYtT5lhZXjI7eexZZTZp6LzKJgoTI3suxdJqsOY5lYObP+9qnCQMqF8nn8pQXjdN
04KDH53x/WuYxDvaA5HqsX70b0RZ1b2u88xZ5vCaE4xxA6rgPX29anbJ/OZeyx7ZPXrLmvCFObQW
A2ZnSC+3eXj2TL/LuQ9IrAB8DqJMbIk5pCvGhmadiR7+mIIahc7mhaihzakBPc47gaSvf9J5aWox
tevT5jbExxJDyPRq0KyQXtaCol19O/yMaILXf3wVOr8G0S7ZuPqoaEpDlQ7YT/tVkT2PpbneFRHH
LsPix7xlymPykmJkAm8pJVrs/xYXx5Zy10uKLj1yyc2V8+SR0/H6TB3jygAOo+aOCCAfmGYZTaD7
yOws6WJT3Ff3wegWFZyvVXA5+rLdV51birhQxHPojebgjMJ7Zs9nRM9hYE2jSV9awD3W3EET6o0l
nPnzKOWyy2r/W8ErHFVDo3TZKTGkK5cMciJBOnLg5JzPF4QdOvsbZo/8dMBQZz5XJ2T5rfgef+a1
bHWL5LfLT+GEB+pNB5o50fRCOdLyldVlp0fuilnqQx0KM6zaMRl6IQI4uryPySXOOZMvx69+kD+W
Vb6mKz8+pIeyp2/ut4LZ1lcHy8GUFf2AN4GU+hlgzKnChaO8Wv/5QP7py1frqI/rJgi0s98g4B6G
Sn6wrVczUkzJH+pFxOKDHCiBImn94thWqtmzpOTWB0pABB/HKcz3zILPt48RBgmbfIvluFI7Fb0I
lcfiYdS8V2vjGAnoxi0c2bclglef1tumrcZFiuOY+H0N1EPjquT7Jb9L05k/Cf1FfXuID6BW5c7V
Ck1X6j7B0f8p7JZD+ieLKPx/99sjnf5C8Btu2RInDINf9TLzQ+Q1/mfHxi7qmRMJ6RbJvT6yAASt
AcOjKwIl05pOF2sUcr+lm8RlVrWe0AVmyIBy35b7fMeM1MTYkpT/omdL9AKeN0eWbmqWeE5fkp7e
QFwbkeXttcU1EB9v1L2qV0UczorwkWSdDF0i5Fxnzk+XbCTTosxcuTDWb3ANh7+FqumnGiWS3tsl
dyencd0fUGbx9smdIMuDmFnJCQHXX9OoAZO8J+Idu93ec873mSrahfRI5kc3TtIFH3sNN9dsg7s0
EP4IGl6J1gMJIkBbOXguBK6z6KMy0bfmOhkPieUr6TcjrbgOwm8GX2h+PiCwzjZ046FKGrzVy/s+
Ti9UUTvifgn6d/NevcZF2W6h8hgIZEpBboOxoHfXXQuKdVIZMaviyssIRLLmbr+wnvGXrobjiJAf
5+3LVH5VXCA5bQ5HnZxgxj4mvP4xcSlj//AJk1ru+nvGx7fG+lQGoX06kPEvVzz4lwO4HvkSJg7r
FAO1TXEtb3+h5ENnEls3L8qfp0nuKs2rPyAPCtpBhxRdUK9O+JgMCuvIwcMpDh5Q2Mx94GVK6tN+
XhamTQnZaoEVWNo7VrvqillloGM+K3hsngTSu8XAwfVFipAlV5srvSIGfG3c2q/eQxY/H7nIYzWE
IVpq8RS1euKf+z0a11I2xL5XpvK0ln+ieIYPq+pr5G1iVN9kZMV6LCdO1/Z4rT3sPfe6/7JeluCG
klRsoBHQBohQaDKq18XmZJGMoB/xzbVQEHy5ymgq1+xS31DjhqpN4UMrP80BqCErcv3t5BmAkgTL
41T1cX6ZZDDJFwsb10J4Dqo4REGe0P7fZgrZY88l7EHZ7sfEXWmiLAkm+iYWUlaBRvkzyXD+Fr61
iYSIqgCfwK4sth7fwtKFoSnezsKAEetLzlCg8cpWLS6SHQZiOiOI241ml9vh3foKGuB5t4auOR5f
MwS/oTqtGh74AkPisHkwkJts4HC+N4kJBx9O04DxX4Zl94ReKOlf9NNdXXGiorRDi7GkXq9ssUUq
aSkPZST09H6HX4NFeqQBeL3gj5loOvxSIihMqBMyhT6zjVvoy11j59P5bTmNTQU2SnEk0PM4sHeB
bgaAJlGFokrbMhclvrIkaLyPGKNHD1kmOLSTSXoa0TATwKI2gNByAZKdFT7A1BltApEThUdC6fzG
AORx+0NKQUXmjxm2rjyKmwXHrbNgRROk1ShIi+58WHcOKCH1oc7mMYfVoJzqqYl7K26+uKmfquuE
R7pK0BdUFnJHAKcmUW1KzMEFSAeJL0Cx9uIH2rWAq9n4vHLb8F6pEi1cV2zkYF0miD6IH3PZJNpb
+qUPehVyOcQnm3eExm9T/I8n9ksM1aXoxZ18XCXzEQ3oncATiWqN9A0FNSOVVcYHHUyUJ0KzEfdU
ryH/WM58ga1lBIGwlyI3EVaadPq9OglF65jZGyRq9e4JBdvs2NTz5N2kP8TN+huzJfDZ4aaOoWaw
KcZyzwHxlEXdXnedqhgJVjsOmAr7+ruwxow6YSJo7pjCDNipdr/Sh4Ai3hcRMKJaQDD+rPHw+p7B
POmcXIHcuLSUtFMgfNX51SXWrTJcSUQUHJTaDjFtqs9gA5RYvuvyMQYTny0GWPVMlbLUOs+7qc+b
hYL/MsEMo97wQ8aCpK7x3FZCkGLnrOTM4kr0fRfjpIUGeeGxySmSS/FAdZSI9jaJkiJSLUIMmB/c
JE7MctHwC0mD3rA/W+9oFxlsnuk3KWw9Px7fVfz150KM7J/UIg6YHRTaCC4sugTn3z8moB/jT/tM
5YrgBl6FBcFHYdx5tDX2waBMPEJJbXZqnJMPlPmLiSpyPi70V+mI2bfOJFmDS6idbswEqHaHUjKw
E1zH7SY8tdZMQzfnRaFHp602XMU4D+C/G5PDFxg8op6exzVEkmFSNS3bF8idR9i3ycrN1jIWfVXM
Pech2tAGT2R7moYWRBSZFqj0t1/R3eYvTUOp1DWSNCR5uWsWqz2E8tOQcifdWriWtF/J2n2Wbtzn
mYsxvZdVkWWq9u+OObGwwRRqJjC8Ik28QR85ksQF52E5uG3ZbfriuxOTJq6SXOdAv8gApSv6hlrl
nh9E42jtejOYE0NHV36SFa8NCzfWRfqL/x4bc4etbc3uL++lo/p9Dw2Nw2VGeuXoEY0RQqYau8AJ
e0JTon1WD24f0Q3qoJlNr2RjDYCw6He35sNRyyWyhJjxqZ+Qi0se55kmB3FzAOvhaqFNjKu84BCs
pGUGMzkuhcFlozk3KOUnOMmKprfSN5uXCs8kEKc7TGmg+aMAB0o3sZb0kqVDYqXE/KS9eFzM9LO8
HRSJIoKP7AkXzWxp9o+akxKEQvL3bgic6WGlF4wpwsgl7OZflK/WsNyuM/JgBwB+o4ndMBILiA7u
JjbgDpBRfE8QcZYAorQQD43Ep0SpQZSboXCIIBwqhFwR9JoZn/hpEMqqE8bgys8uIcU3QC2BOe76
tBH4tNCu7JY2OVGnHhS9Q1CTs6IIgQyPaNCHHGhIsGyvxTHZKSAvBdkYjxGRdC0tXg1XXPgRBiEx
/vG6tKL5Wh0XTVnEKfwYTeLK+dJMptd+NlntxEFQkOajaBulcDkV+nSEhrC5RNOzCOT6Y77z6N6O
RJCew44Wqnpa+wmiZzBD1h6lQYv1KKJA4echZxrrV+UQYruwKl0pnpew4jwlRL3B/q13pfuGGKUq
3MWBgRONxaSuOiRSHI41YztsssdrhTmtw2VnTVQ4XrpF0qIYdooCHfzDu1mudV1RIsOY48VyB8/H
ghnuoAwUWTTnXxSjLQH/IsYINZFDH/RIUpzEolf4OMJAgFNX+DF+oAZE1zx6MROjLqhewQvFo19q
PpBrS3jURraQVMGIksGOE5HoeIOH7B321dfk2W6Y2eg4OugOYdPYOQXFEmM6z5EFYAjwrOQYdNUt
5wRnpohfwsOw8ProKZsdDTUvKurM+4sbAwgOP+cS40+10PgvGvQeF4yFO25p9bnpW3NXlzhIA82d
TeWxoahMDMjcsgCB2RM3ICP2VwG9KB4bMXvvJH29v2qXc9o4Zi8KbAiW7GmQ/L/dRu3hhCdfhH1p
YG1NWvlRSJoEMLveDe7taS1K0eRkUpTC+FrDNvx3NL83GXuCEEwYoZeyZ+rH+Aim7aVNCBaPmOS5
C/wcVPNNHIYLwcWPNNpgoNEzUMl3BrLX+dWD+WSMM01WeTdP+VNOuZDYpG0rW4gurjWMjUk8okAH
WMdhVCsBs8WzEd5EB82+WBBgCxyygI6r3Rf2CZbHarGXKWgvTPmbF0GLUEV3VSR5fXvQlFSr+bNt
kYPV91IiLJ/PTm0GHgjYut2Ajgl+Zks5IcVFs3i5BCEx+inS2v25MyMZFhWj1rhBVy8dudGwqBuY
9bGGZPmj+w8rUxWhxXdGFdAyJbf4THhDKZedFrWWbJhWyRi88wZPdu4q5ic1q9aTKpZajStpqMwI
LGFQHRBScak6nq9zqXS/0PcGXMnmNfCNnfwN7yStN0hFcpp62B412ssSoHD3O1GxUIkBtHwBTjhy
LI6cYKEGkCO1ibpJa+/OYrrVjyBNX9dHuWLgp/uHbBg5AGUogYW6hDXChMT1GCdx0ZJkfUF9mF1b
O3SjT6DZzA3d2uo1B5XMmkOTsXjyl81FGrT9DOf12pLcJHbH6HzBytv8noBGNRU07Bnl8eV+LiDS
SF4A8UF05pFw9ZxlPuIRwLjQDP8FqwWNo/gOlhEPYAhrQ4Q0qC/+5LuUe/0J2f1ApCmG6N4Kc5w/
FpDgzeJbSBmjrL0x9Y1LVQbEpC446i08OpShl9IALo2e04zsHTxDw8fqqW9Zwbso3GJX+wSL5TNX
oB8MACAlrAEyWHFbeJteLrhHc/FRRj4jdfyb6YuODKCNiHKC/obs2sI1FHTX2NGVL91+GuMWG7Bn
oj60zz1aohOY2LZr+Mntr9lYN+MrFDVBiugI4CoCeQB0ApYMTns3k7BRvk6tTMVQpsT9yZJAyRBL
HgyfLm/TtAPMyZdilDWgpcRWHU6XlfTqJtO3E0gz0ke9vujlJCmBT7/1uZ7pBXRBLQgj51C1WwIT
hyNAXNeIbMKn7YTYfDNT5eV0VvCKXW9bQdsHSndPPEgSJn55SLRbvjZBlQ91T7xR5TOUhJMZHjRU
lwE0KdhD4+IJgVZZCi91oKzfpm117doRWVfWDa5Q3ptal18DGxtIZJq4te5pQ/qPvQw6uySa7NIW
rmLvbSUjpZ/iGit5n/fHf4m/im2vJaNPPdlWXDLMKj13bS5/iQXAJgflcM3xEDo2uIshBxS9lR1o
Cn2mUQJvawgHqQqWRNXUFNkztnEsDIRO1XqcQQPpxB6COpaywodfAdVHo5o06JKstdubMkNT6+IV
fbt6lpylOHdLZeNpU4ZpzM34cENvLYlk2tdrp/KOCyHELokRmmcNfvhMe4nj6k8L08oKGCsfl+xZ
qqFNV0nKuaAgUafSpNBDA2n0DeTzxp40Y6zyAWree77b+R2VlNW8CgG+qz5sXqkpFLgDDGnuCd2t
Ixvi6st9cAwP0Zj3y1rlKgUNf02BYXO23y0btrKeSgiYRfAmnWG3Jn58k9gQvWEeH1BH5sgrT/Xm
NDH73RBSGywNpQE++RYh/4zR1pgE9Qtjl0YcUt6FqQR7sj/BEuwVzJSQRqsHIvk4Fuei6WMGgFe2
wO2c2zxRdsEUkLaPeVnV8Rk/fBfeeAqhcwr1KvKvPKoPCMfXiYnc1XH8S7KHzxnNGVPlYfLdOHtq
CjszSYDfE/iYUzu2M+AHzQZlwBVSIg3C35c3SCJCkNH/4392HsKwF/wVzEPi2wwoRMWoa553QuJT
0t+wPJOkOySwk816I0N3a/7bwikVaXTtl20girh8hr1jlh5jo6cHumOYZ+J8VFXhGzVdEABNnhHE
54gY1q6xBJ28FN6kSrHBROoGPRGMtgeOTqyJbxdwwME863TuV8n2FZVphutfBB5cC568gm3Vb/9C
MqQqttO2wsO4YqcjysmoRI67te/3/4w8UjGfQkDB8SqtQvMYNj6r3yctBaon3XqTWowWPpoBmpu9
qMNoSVyb2GBGxyc2fGTwUpYJEE7GbrK3t7F6HJjkV67Wv8uGdhN4SSTlzczKS61LNFUFhUjCdmKV
6VGwtstFSQAla3+tgbUhItKfWhSHjUzDYNg3Tm0zEOc42ualVEolOTL1ZyNp7h3/UiGgJXs09wLL
soNzetUaLZkRUelXDzgx+nNYLPJxPLzgWgBAg5NhaccycisfYbD9XNZUMMeuvSNWU2aAtsLIM9rR
MNnicFUKkyE1irys09qERrrWXG05ESiDXFN1LxwDe/D9txK9gBf+AECwdQx2e/qnCONiZWuldWjs
Qhc4ncqhq6dIvfcMCijW6TQdx70cM44MIfKWrxUDQ9ESDzOcpjygDaZXBAonWa+x0CI5xWfC+P3C
dfHZ6ENx7/obdXUB9VnDSZuNvDBYKr9qHNCWcXxQD1M6mqb+m606NlZpeyapQH1897aZSEiX7DMK
bFFzSvhSfBvWqVUTjguStgAydkOhp8yPII9y/qOQvgoRt3uldIEwjZmeFzeYsDwp3Sqz5H9SNXtJ
RejYqiLKjzrhaeM7E2GuCevsZ1gCI42Z9QBLmK/ZZ0X0WmU9XRWNV5k/nIZA5Zid2nlCKrn23hDp
3KcImjJxH8w/PcUnSlAPbzB9VwG5YY+oXeu/NTxyPRdBCYUPdywL0JPpDzE57C6s1o5ZOFVFXTtq
TKf6vzSwRNEmZusB6phNxa2eU7fQR/+Vo1fRvJIDY5D5M3TDH3bteHAL8hXy41MUvV9Jcch68YZN
7zJxFsAQ45Uv2s86KdmXEHxOscOAqEjvM2qhNWtrn7aWvhuTGvOmRkTN5YSuAuQ84iIZ2JndjkY1
kNur5ksJQQZb5H9SDdeCTu68z19r294vrQCDDLmnLwsXApoWiAFAulzewfa1QIlQIG1AkZzyUP90
FbDTZvvM9Hrc68N8kk/On4WDm+3Hxwe9wJL0ZldOKLCOEpqTdfkyzeZSBqfprn0lxcKse+BBOJu+
pp2Y08C7uSFnlFQ8b6pt4wIRIPwHScvVH03V8CcqXYmksUAjUdyhccaPSkK2iLtQzlij4eB0lvc1
48FqF91iMA6MY2sZnQSkCU7rL1KwDhTsdBZ5vEmpYnUKDXJBPi5dMYl4iezHlkKm4XBE0JSySuQb
OhA1r5Dv0fSzSekx0ywSSeNSsrBpfKlv3EOZ3PE3wb7AbLgLCnm0NE9nYuuEaWvOWc32C8nKtLTU
MKbyxIXMwWRXZS9oCYyp39svTiXHVvtptLCiScEkllC/0OAUKKWJPtv4YqkAWDI22J7I3dhWy/EP
iXUGGdiFR6NbC6cEEbBDSD+SqcVHudyYB4JWrcemDRSfIHoJivRd1cdZ5vCbh4hPgeHpDAgmsIO5
Scgkq3d3sjxn1G3J0t7SezfRKea5iASjvfH1APZsD4MjuyGEYvfX8gJeX1wVa4XeOasgfirgPfS5
WpkYMTtK4Hd8rQH6HW1H189QLZPMmU8Wv7uxsYS1AeMEYCWw1Wwa/7Vk+9xiYgGY/q5Edx0UKG27
5A2gFqxXQoUnvRQOD+66FiTBCF4Mxw/FXHebOdsK1c+GOD6CRbah/BpZkuM1vicCj0A2N5YmR7/P
OQy2dcOsrphrw61Szx2APQhf88hwrREzzLL9p3eVjuUxhI9oogtAZzxJPtFAQL+slyh20Z1aBIp7
Vf87TPTZJ9tFXT7z8egD3pvZR48+Vcw+OqODfMTz8Aw7tT1Owpg3FwW/cO8pOrEGf5ubuRKgvNI/
u0d4lWm/GuSBj2ibtgP5+ANa39rMLD5ty1GkWqjUPU0eJUQCLEz7RU6RcANyqEsR6gFVDwbXeLeP
2r5KWSuILStdb2nixaQBnyc9EOk4Zbt5HtO2woKGlEVxt6C0U51hbExhWl14Jo/gXSEzkF40hca0
H6Rw5Ictwp56LvjbYHrIry5GZTAwy83dMYuOaCwboIHZCASGj6PL5xbgQWN4p1Gk+U4RDuM+iZaN
+mv8BnGY1lQmo0TvsNTs2touslCfQ2rHfLTXHTnYhtJimLtRoC/ro+JeMERMNOksmwLYsYs0OkUI
j6IIqjSnQ/T1q0xKUEfwtN7EuvHi9E/LRgSx15YXPGJ9/7HYk0lbCtPVTW8YN32otERp6rmWIbTv
nhTbFD0gWklGrNdhkLrfbf/oDRUoyhBELzDx441NsuL1HrfS2UK9NB+5G4m3w7zJQ2haJiLArq9M
lYtD9R7y01B7zsIhNhGxbyi/sVZP7gXcEmT2Ia4QU8CGJUvCxN2956tk6hMhGG4IXf3eRkO8lP77
1rWP3npNuW3JpDZ4jyeFuaL0CXXxrvzZXKVMbBm99CLCf+FWG6fyid8nOarEKfn5yNZfzJoyQsD4
nE4mW6Of+i7dtZF4LXNcdgCjnZ3LOt/R/YyKgEY4p55VuSAXAzJKD0bHyQ4GIMaSc6ZIwzenxg+T
B2kUWVp8KDf0uc1zoPBGtszvKVz1BDRggE7fGzHAiY1zpGhK3krGm/+vhQx4+cngrBax9YLZ40Ea
np+9DZjh4jdIAOYqlyGT8NbfGfBYs/swu83b/aYXZjPYT5xhM001Bk7j13iK7Zbep8jnDXRyJLaM
SU4tXzVdDgHOa3TuG4g6wJJqljXD0Kg4ISGyPyiLk2QfdvF3C5XEz7pMYcpd24qwMBYnwER2xzp8
/GjLwkLbTKoAvPAFU9ZDyGiiTwLYkyBSLpUw/wPM5w0ub0E6G6iD02a+d56hXejAFvWIjInHgHED
55nq/9/HYULuuINOGOhZr9hF46fDsta/HSGB+OjFpjKgCsAGZFTFg+fHBt329u8ZDcl2vtYfhb16
oEcHioP41WV7kklBRDXDEuGwCtZ2n9pLWII0cu2G31uI40v6vi8N+jhIXZ1yGrDbZO4MEUUAqF0r
SR+EbocEKwsz7EiT+jGLZ64UCqeVA8YDKQG/PElb7LhXGhK8SlJVCsPnuqLVe39SHC9s5fVjqjlZ
NH2+Hz0xGRRelCC5og/jec3gZT+bJcg7AFaRTRpQup7T5BATlhj5Ur9Ulws4FktpnIvywFirCgDI
UikTBubq0BRiifgaWPioTWpBzqlB+VyxenUZp9C50lCrLfxf9oH+0GwCnoVZ7C0tZs9v6VpsVFPb
9L01gYnLRfNEpP1ehPrX0Jih+QsbR1NyFBgV++fHV/1TB3j6As5pgt4uchHxcbwawQR+60loXHWA
/w8vkgXk6gayoQ4vybKCZ0guWsjCNrcVv4J6bMbjsxE4tmzqK+9cvsu6SSC7nS5Gkq9ggSJeHnSr
+a9b2oH4hw+9ZpzVfWnWyXcCY0Kvc/4D20Zh3eBG5Y7IS9RrI4oAz6IHRPWu0QUbpB1rOBj3np+k
Ru/xnIr3P8jyIrDmHxGn1ii9utawa0urioSnBUKOZlUtmyo2kV0xb3TkWysVOSt/1x6ndgGkE+Jf
fT7j3mZdOZN0nvZND0mx+M1Z0+W2kIcsQfVYB94HPNIh5nS80LQFkSprzBjhGlhXkVNkrHP/o8/N
v4YvMKYIhlNulBoFCDzP9j/f2Lfizi6os4ltbx+m/rqYNmp0Po/NWYooG4BlKbNze7swFvi3o/lY
kMlPpWV2JoW7sPZV3ATz08tthRQJoIdNWxBZTnjJu/4Qyu1/8Vnzo8As7uuhVcSTVRmGgWTHv1yb
jUBnKkiwLu6CNggJ4+GwGsBeHePNxYAFj5eBxC/AENPxp7bA1pKUdSCxXXqYtkxXhwO2nwG0TkGI
45ESYFdw2ZyfVr5VGz03yzLKVlJGmCJWudKVvt6f+NvmorxJ3pv6z2kfe758OJNnvw6fNJt41UsH
bBhhYLNC6R7jj1MkyuE4oFPIBn2ba3x7KuE/GYQj75T28KL3fS8J9kDVt2NdrzHMODC/fiomzck4
QkH+Wd/gQeJBZMOBi7VZCTwbW9353fQhQ00X/4RYD9UtQZM3+AcaUVOAFj7l7D8c+6IBsQwOj3Sj
zWi/8TGl5L/8IAjoUC14YcB+2ZNdj0+EWMNqQjDxTKAzqqhNG8SYnFAHby6RZdUCJ70vSy+p3yle
yp9oi4/FM36tV5DjExwe+fFBVY1CBBt235Q4BScb6oFd//M4/tmu6lrhepyWjxDG44nutXjvKJ8P
JQaVnEEjsCIzOGve+oLHQpWWNdVfHxvx3YcRSQGyBWtLM8BDEpsAw3Rl4efnls1XP5Q/7M9P2q3/
U2qfdzLVc9kyhK541vheIsYOjJdXOSIcthXHC+ebpAPCqENEU6k3maDl//Wly/8XlaneCvBmT8h5
12u5ejKDsTh/ZC5PogH8xtjogndXF46myFnEeL4TqsQsO3yUbocaQouzOkke9kg2RwgH2TOsy0wn
AYVtRv+JhA+uyGkKv0O3LCRDQ+sWBqluA170QTv25Ouo7x7CqdbwLjpxoX74t7wJQbNSw1PhVQze
iq/mVTBbe439r3Z9TId6NQtOaJ6R7hLY/xhZIRx0Oh70/PDVah8pYqaEM3X3Ye2IcTi1obpWnS3m
XpBLZ7oLdxco2GvQjOAnZftqtk+Z+PLfts+M9si1Jr810Sec9sEbVcPZTIfYQU+Ax+GKYcOg7HXN
I+Pucqq9vO9R1HS/YzCoI1qrfmkgKrcJ8aFOFaqqTDAMJaOlL8e5CfpfAWqFjEI2c/jDMMEJO7K8
6AG6AbEJ4iyA9U3YIvilvY0DHrInSXVpRpj3RF7ughaAHXZrP0F/v59M0bqTayuUlbF598ojOrj6
OhoqYFTw0rrUJLj4+VD+rl4tMmKId1UU8IZlYUkloERO6D9XKUkaF15weAeni5ZelMMcspXHhRy5
XtUAvAB8xiNoMKRKQqxJSUWu+UrQTB7gB4kM9UaS7YFToBBjjForvQBCOOpX5UJAM0jc8e2egl9o
8N7Cy+Xbv+BW9wkanhc3rmJvdG3xMJPY19r7oZ0b0xIP0WOa7O9SR9yhdcHf0y9p8L4HmVsCidBx
EWxckfNN456mX2UZr6+P7dt4TCHtniu8HGSh4cCj15/4ALdGtkTFdhXJZtdY/ocSXLKJiIMIENnG
3/eVyk5IBtmagqFPhDd/5D9EjpL6Gy+5sN5RlTLV7C7J3eF3VolZte/7R1nkYCzpQmmoC4q8pfQX
abcu1nmUyNiIIMCib/ibOY/j7jvSfAIZ3HKHtmBB7fDh7nVU0VkYsaTk2uL7m1hsWgUYJMnju9wG
5AeirgCXsY81CLLEoYFaOjY4LXHzgzojuqyY9W0AlhYL7QtIjsAe4AHghmTNzqbo6BYJkj7oZaog
vHwnMWarDtvpHL6sKAEqJzfVe4nDBepcezk0OdCs07xU60CbpzrWquU41ryY29qQDRxW5roukvoP
9/RmQrpk0u0dAmGGH/8DurJ6F20ZJ6M4EdiZjpLnZcAohKGqqp81OSI5m6OPpi/F7GJa79S6VJxc
nOuPv5W/qUmfWqO8ZV93JmXBfM+RjADVdJUMSBnIicFzXhzNjvrXp5UM0Z+gZp9it7xmc7mrveIK
JhD4BbqIXAZAS6ZzAqJztAVA7FEznDtJig+xuwDXPMQw+Wcb2O7ST2MKK0mnJwzznEo6uSG/iKpU
8Uo3ERN2NDCvpeVx1Jbkk71I3Po8bFnjlguJBqKE2IFprYk4WcL4fL1raby9cFSCKPUxKr6r1b8W
gCjg0ouM4nLkQLmkLcTWEcOeizN0vy2ROaE1LORd0e4bJKjSJiSlSlyub1HzzovK8SeuiTArqjP3
jQZ0Psn84sKhNHNAzr63xMynpYmZIe19PG+1nlIVMAlLgCGFxYElS1nC8cwiSghvRbjzd0XB93yW
oodCZObYmv2XJ3LDezU8ucvtRbTzMxolMS+jM1fbqSD1IIw8dgc/G2191o1AD6N0YELYykhX6CYb
h/QgT1zvrA9lcecCIx3VaIbO1Yp8HFARIeNhnJLaKXAsQ0nh+VAJWEnWKYkC+s5sGZkGUzzOteUA
q4aIW8qbWKfUXEECgUiqv3D2R4H0QSMPcRtrc9/WqZe4ukG4hJH6znlGqUAqrMXOqrqeSxhWjkUM
8s8U0ODLsoj4LPeLgWIbWhDzx5GUfG/ni9Rp8pXngQFnu7jiUIHJs54OHXy5oxHjansq6+Pyd8c1
u48pXbTRgZ7O6sP7xMmQ1pL58imKv+6MK/0sLWzvwjHC0N673jqpA5BzxH2vRF3d5KzYDobVO51N
inLgxoU0H4pbaWh5N7NSy0GMRAQqNccyPTFLmDgMyg2040UyJUOCsroUWovF4YEgyYp42FR4GT8F
8q1a4/KXie2IxLdDqKBF9tSQJ4ac6Xs290lQbMLXcZlMzo5Oxt7l44bQhG6WObdCu7OWrPk7iOWY
TfyCrFEJojnr4/5YTWtxbmLjPXkUbp78elLDRs2qD76c/jzl1Jy1ydhVhTWfZ6V8x1QfMXj9L2rJ
w6ueXH33AlxMzIqX62sZNvXSZhaf3+3hJtHfXrop6YGC9R4OjXdVfVQ10AoiK6IUMxgkyTV90Jnl
a1fLL3hIVl3kh8mlf4abt/JWZNcoQKTO4bzBg3u5R37JEtUsniMmk9zvqJ5PJWI5qBOmbGwu1CyC
IXI9rJH61vm9iByIAFBTVvu7MQ4F+xY5i2BZUihyIPq0RUUXZ26R5EUALBADt/8/VvpOyjT+JyzI
Qy094IfeW4GGLWkeenU0cI9XGTUH24RNZ/LwkiIw+WBwPVN5HqC/kOCy2/P+C3yFh1WEWhJxg1KP
Lg2lswZmRt4BXELtb91gJmOSl1rgHEv4mBPefxdfpoJhuqBCe3jAt1RMjgj9SIsJ4tukIPEyJ8gQ
OT0/fVTs/985KReALPW2BbxO6EBfbnjT/UyqprPi+0s0q+3GSZIefk0ONnPEelWgjdPbYBRtFhN9
LpuKzSxVkhcuhnzydOr74g3q384AQVC/aDMtafyVUhHSxF1DGSITt3fY0if94+b3OFirwAwFQeZK
SfefU5bhll4HmKZ/xqHwGjN5rCzBemtOG/AhBohMT8Hhj8a99EZ7WIB4FNMtKwQ5yfa9Pd/o8QGX
M7+B7pP27LUw86WzolCI6pQNsPCdsNSLf/hx66K3BdFwqWx8qL9MI0jubNj5YBorEV784N4C6xet
uJuXFvyygcleFxq7FKtMUGzUUgZrYELiueZshhgTs4voMuXhSUXRo5kgTg5atPu1XBWDKf12T9sz
/BcTKiLKVIseVtfvmth3JoA0lKjOFEfIpDZaBjF/yv335t5CDOMQ2yKBjpsHKIH9x+PPbmUDy8RM
XNEecBXQ8XVJQ9TsRiRGMjWtSPahAcBvS3m5aKnvMn2FbbnpPmx3w56ukeFchG0/1qGwUyR+1gfJ
yMeSA3z1huajEwXHiSrtTlCSPB4P8e2jCovOF80gR3adbBcJrWZW8VropgabZMth9LwS906L+mDZ
7q4Y/NghTfThIxf9m4yFQUD5RaRWhBW2F867m8ug4ClxIyN8R5Egftz983UdB32BZzObmb/eb+w0
TDXTZokFZwCln8iFVUaECMf0O8gPW1Oru7y7nejDt4lkwCdx5vqXcpoScsVZIGTszvBUa+ElNMIy
FofkZIvLxw74susPLfV5GLTnbA2XoprFwDaZcGzN4glvE2n+0NDLLX4JBRrFaSejekD9abrBceCO
4LUtTFzwtDJ+uWS2BgxQKda5nivG4a7v342VDvaW8FRUWh+fGnkVFwTLDZigrUIquU14JO+cmhF0
iRKppPdY565tKlY3DTHdeXts7s4alIGI6fijvzNArAtQDyughofcmzVEFr+fXAsnrLW5kH8IASTt
Kk7q34gf/8RDF5w+DHHGAMftUX46gkQMhYaR+f2Mm2VLFUbWtbZNqhJ86EZuB9qpoH9cQvWwDOXQ
UEMZOF6c8XSUh8Rz0xCIKRS+8g5J10yb+9gCysDXZRQrn+ZWk1ylz9f2zBpMJGU/xgt1GTndF7rD
qGun5JKH0ptNQuvXA1CHgXpz/DxYzExQ2uI7pECdgMWqkOUQAQxt5VUMEjmjRpyJX6/Bl2TtaMyo
k7et0OIgSlnG1Daq7QDrjKM+sDW0KIoBorIDeaN98wmKO1effinT/FUGkY+fRnU3RoQdy+SR3iLX
1thDxfK8MgwX/dW35pElCzkApTN1CPCwetxre9klOLXeXdcntqaUCWJ8XPi+iy4QG0VFR12RoSAH
sFJ4tTbc1wwoekFRKGOybuEEnfi+7WVCv+VtynoX80SuvF3PQqaX/VGDTbhqa9wFU7MChZpZ2VkP
vPmNPzj+nv6XUh8gvVEYgfRLDSuR+Oe2tZ6oRw7tHNAKq3GY/2RY6yMcPZcEOICBWSinhCjnL00z
IMwIVCjedAToral7n5Ifx6c5m6tOgy99XKBr2WFSPkRP/hWYmuo4s/px7Aj/f4mhGrzMISA2nQhm
CtZsWox8aeWKdsGAKfqI2CfxtPF7+ISREU6t40qAP8S+BdOB0dGxjcXwPVNtvh5Rck6PkiJxtZn3
7Scxc2FtY2HI9esuJuUyzsOZkS+mi/1P200Bj4psO3Dj+NTi6TXYxOuTFVlmyOc698Ys3TjB0+J+
WOq2v1IQWVHDYX001Yo4EzUatil8uzJmiiA2qf4JXOG13RqodNnmk5r4Yfm5H1YcMN+TijlKG+mQ
WEA9cOchFhbOmIMNo1S+XIa9MaQ/9RY47/978FqY3d8joOYLydiqjC7OVm26z548+pAG0Fkh8Jrl
1qcqtY0iRusSZL4shc4YdF3l5y7c/bZlWN4g+FSGjbgXQP8SwMUc1tSdi2gtKH0Ipq95lOUvDxYL
NE4V1vyZbBvY5tKcO1dByUM5WBgiZLiWtYzBfQ9A8rISozb9QQL+AfOAWvvgCiW+ezOTLmGHp+/r
3Brc5R3IKqMsO2bumPjKRWUsWY5V797rkNXJ2SV8x2m+x2R9Btivf3xBIrBOMuF+RGrujSZ6+JmT
NbhYwCV9G/lr85ACMvL7qsd8aO/xjiU5BhlOGXZM7D9hHDumu4Z+vjc8orEY9kHbnyBwWBmEN4W1
qY1nx3gDQwsdh+KnwVTgFvctruoyH0WOLDznBJuGdsdqUbZqWlRORiqZJWNCWrMf37zA1HfrGmZI
GtU5RkVSiJpdHfciwTVzrx6sRY7yMndP8zLPXDVXJ74kUn1h52d9gKm+V/WxIjZ31lkiK5c2xSZ/
tX6PMXh6MPO6CacOWmkYl1SZvYbk35NJK2hC7gKeLK21eCNVE4PBawj2D795E2xWI7cgrdJ55o1P
AfgPSSUMoWseof2ikXqCdiLXDa05X7qKsiYfBwkqEvqG6XrUCdFRqGAWZd6aW/13biZFL1RaEs3o
VNqO8t4TI6cPQI3XRiH+pLREXdQTAEM/yYg+XSxQxswDBUsG9Zvy6gYaD0BFmqsdGDWw1J0eKznJ
cCXLNGFytW5FTuc5xfHkGZzxiCyjSJEgtwOzP4rv90YiGJtOp4ZjV2S8SA+vtbGgV5i4AIYDoEXV
OiIrQ/HdA7BWdyNWSgW1VmWx7emZ61muxj3f4+jKNDmB74XQLHGRLmGD7XFWIhXEYSaXDyMu59p/
heHn7m5EUpYEAnzltXeA6CGuPtYjmA7dLgZmuQw6qY9beaqmtUEXIaq4KY7Ume9l3SHGQ7jxkuIp
JKBe1l4slRNTZhpfKlADsI5OCYP/Z5kLF2m18LuVcfniIwQkdZJxq0KNdhKxdK/vu1UsjnPm0/6l
FVAUQR3FTMGVPRSYTXmfxV4xqXSi3CtCxVtWVl3JZ39ejoCCwL1Kd4sDflEhoe8lzy+4YUhe3SaH
v9n0Bcx8ykjX6kdN/UMjGNW7N1xJhWTjTDO3qccT3A2dGUV5oIyjZFd80mRHW5Xk7WdW2+g2Wq5o
qNFC712olGJNTRfNNacNcHWe5nUQgaTVxAtVDPlWH7yshcU5+vRpX/E92h4h+H23uEZaZnkGS2HP
imIEeDOq5w1GTqNDG2agIhKpoQWJgzHlewSpflDHOIYd+ANC7iAaO5nBWNQQBuvP0dk03f21AJmG
oqlowIs5TJiHNQJx6clIRU70SXUlwMG4ETmKIAq1qzhgyqaCTMX1TpEySFrj+WGnOOLTld3+S9ps
eOBhDOMCFLb3txvVuDKrNMs09Ggyl4FIKXbQ/7eOVFBgPXS96q8HtKdPcqiUMsg3uzJCXKX+9o1R
eto0B4Zevwjvl8nw8Ow0bxUjwrIzhA0cHLqhzQ8QsojvJj26ZoAeembpNMRAhbtupG4qmS56hiHj
Rzvq9EVsevLPrDOSxnxRGkKbEZ9o1iR04D4zBryP9Z9w+gUapDMAjbw8j/eOOc6MjgXBOt1zNWjd
YlkWeEcApRcSthQtIja83br//bu28gqPigizU0Zas170Dx1UKtPmpSB1YERhSE8rHyFXOajVYqvo
J5Pa1yl7ILOIDfZF7uIfYjVa3hi7DxcxUwPkdYKTIgZhjSwHlKOTbMs0V4FVKMe1Zp8DbnSrwq0r
LX8v4s/XtLKRkXEc+IED+rhSbw3N0p0WGYCs/+56o7iUtb86N/dT7E/d9IQDjSV2QgwnFiusIxJL
65gUwtOgNdWMYR6vuB3RTTjFlqXyshOgdar7pf/Tb5ZWNsYvZ+wKl/oW6kO+3KJ0lCBEYahZ02rr
dMUdhwPkvaI7PEqyb6nh/dUHfRq5OOhpRiWUYb1WZ5tLGuNDHIlGqCR2A21S+WHTPs+PKftN+kFA
8msUH02FdrCGLZjRhy+dA0xrYUALkSseqJnwNWdtGX7D11fYtwUXE5cl6KxX2WGOG4c5+Faf5vw9
HPbc4D/Vwd6OC+w4cQpWwZ6XqLI8lesyUaFt1D58Ow3di2ujnRPo509dWzWtrIiyW6MNZTKmj3NU
YXZd6uMPyWBfrvYx1AiipboQimL78KeMJd2HLWsNzKerIhyutlSmJrPsh4ZiipWBtXGYQ8RgW7A8
aL563bKyQdnVFsaVQ28CJ3m955y2naLys+13O6XaJNXRSoKG6oJ9ZbgwpUCLA8h3/9NlmipThJP5
tyaLKmSJfKJKEKMbBzIpxxeuVzBA3Z9Q1M9/8LMOjcKLXZ8iZjrikoOFwR2RU5ddAzmv4svzkbOi
Qo2yTMetEjecJwjMGJqr/xH8f2bDo5gk1FoDFb5PTRU6sVP14U4wnmxhP+sE7jPR/KlSje3l+8F5
qlbNFljC3eC8a3M5goolxTMXvm72gAk+84frKaWQSMtzUP4gyt2WaqKsVBsOf98eGDxgUVUm4TaQ
dzgCFQAPO7j+LHTkz648l/6k4j/umVk7aKQT/jdD++JopEvNDXE7T/cYiUOOhnyt3ph1KlXGtHsp
oo6dEEXWtVeeM9aeDDaECY9vQKppCzZrYSBi3eaFhxyAQIUboyZLl5S/9sCGDh7nvCtLHjj15Wee
y9ZSUG7X6GSDFj1NAyKsvK0sOZpSvQa99ICv53kOFEgPbCjNguuRXxVj2TWxdKNIdTmbXDD2RzjV
ILclx1taUig1axyAPlm7VsP/AIDHf9puok4q2zZGVYhuzLe70cv1wBE3GFbOV1CDkV7UZiok8iie
03AZd63WtcucbzxXVZAZHKob5M+6aSDJSCDp5BmXmlLb1gjT2uVYoMZz/c03Vm/fh0cwwnXj9FKp
swl61yOpks26Nxx2UVhKVE4STbm75eaA+ZnHROttI70zhYtrvecaBDqOI5J1nD6FKPYdwqXeHRky
MFryYrSCilPwxG6pYaShnBj4eyzsonff8Zja6ELbHbCf9Emn+/JElO/OnCYQiH7aHoI/vVLYGgZV
GoQuKBxi/lfh4QOtme8fdhiJv0rddyd72WkOAO9Jk02fRViVu4tn2skcujjCIi8/McZsVtZKZENK
JMj19eV/XOmlaii/GZOtUEExoWoDnSR1BCxDtQ1Q2PfZ68LXEiNB4IyFJdFNzZUbIh3tqdZBrtWS
A0w34Zp2jJiuiPCNGlBbTjwiDBsJ2zW298ve1MmhOQX8UAipnS8dbEvrKx8pp11C3dA2DmW9+/tu
CkhCVTHHbZ5HBwhO2v1DT6JZKH2KF55H1i8CTlcGd5gJc7Dzc+3Z/giWy04LYI1uyos08KY+YjtI
R5rWgRyg6Mt07JUH5nlIjV5k0n8Bl0E8FDmhiz7PcHdGbIzzxxGHMXr0sYI1Sjsh50nd54HwJwLr
V/THJuXcDXPqquxwxF7VtHE3k0Swl1QQBqG2ZrInWh8FFZZxopv5T2bvoVrFhUHJstfcYdOY9Tpx
mmq7ja7EJy9WqV3E900iSrzte90mtJ2RjA+YJk7ofU+Hrnzo4drUa2ETGZsmxvcT7mEY7xrmC5T2
/Zy3QSor+kSVx900/BXCwll1PoBv7KYqobzug7M9bPrnp3OfKSflnr9FVm7Rr3E5ao029CATiDiE
6rgBjD+Sd6UzJeBojnslYOTNTSlOjOXFK0+oby7+4BwFaBrPvqGdsNra/vj9wKchX5OoKiXf7wMd
+f2paa2KWS1BPGKvbXCM7ne9nsqcHrR7Rdq8XKJs424XZbQl6Kfe5TxZl4P7hv/8d8Dy7OVUoHC0
OgufG18f0Lz9w/IkYDKux3xpJkJJAzHuR4DzCdD02CAGiaQYL64IRmQldZvmWgt2pjEPZC7IYBqI
XTgdua1Ys5xdTroz4MNX2W8kdICC1Tg2Qsysr5oZKSH6mqhlSjhsIGB+qolu8a56kTrXL8HMMcmw
6OR63yDTwDpxGrVtiLm8p+F2fd4Oe6kbejnJWZGXNU/IP4mxL/6wwlD0pBd0UqQOHwJ+VK5AWaYy
YA0zDJS/D5eLw5adODOA4W6tpqIGYB1kJDb9fs8ZEUCtpFVSxKZxiq0ViqjYbqrIwpp4Owumo67Z
HNxbkiHr+KZkkGcW/P9yrKm7+dcTBSEBFjfP8+sRdGpU0SvCV4mkR2NML51Us64BkyeroJLyl2m9
GJvK1PpLuzgeJ9hl8vlCufY/VkrDGI4q1c/YfM85ApylNZ7zXiDT5nkpLB0Ga9p752vkvww+VYE2
Z429owbHz7cvB+mRD/W0YyHgoBwxDOZMaIQCKZOuHfarrli2Lu9ByvSfd3bp2MWtKGacj3AsJz5C
PP1x/0M4JBZx9xNpoxmog42Ju77f263Z1L1HGyaZSEZaaLo/GJJsN7a4bgVOVLXKlQIva11e95IT
kSmfzgoWFeUGB7n1HAzwpw37+Rk/aB3CVi9UJycCVtc2k9elcppbyrru8aC4FhbeQ/mDJouPr6kP
tyt38DKMrQADQAqEfg7f3oiOql5WmlPaxwzDuns3GBSCvNWqng0bxU+M0YSBm1lC8F0kBmzFJgnN
ALB8J4uTYFMjhjuF8tZFMJo/RYQk4Vq85eVLRYWioRvqOgNQ8z1loo3ENuBLeGuKbaELgBKuSGiA
rkSEueqIMA2k0YCfE5F9auOzCJSiVzrQEXNTAWe4u68fWvRADz2YQgX2JVWibhf6UlyuqurgvZ23
l4CgXg3tbTxRmNS21NJwHmflz6pPXp+TvVVDcVzXHUJnvANnPagMSCuNbTqqxKF/K6shjUW0ebmj
+Reln/sYSwge399VrAG38iRpOPTsB1ZBdsrid02+CEGI/BMhMdFlp6aF7GLJGiNEKBx2D17BjCgy
aO7HJD35N61XlwFYZW1rN6uUM7/FligH+H+2lou5yc5drCsKjs1r1WH3o1LIp9cwkdbHqxNvK3KH
9FTzHWj0L2auSQoKDUqgGsz3QGdsyu2fGCwF2wL4H4VHGeTurQ6h3kOcwR40Ys0QzfxTQ5clDNjo
V2wGe5E43uVh9rhXJ0L8goRp32LSR8OYVd18OTMCzHW9qqjtu9C+B4inoePOU9IYy5zRGLLgpS/b
ihn9DVLhyxIuZukoj4/EvqThXih8gvDBhzhhbXpzO3Uu+Q0LbScehRACeUuAj7G1roQ89FbSsriW
gxngg08A+Ia8JVA+p4oMVIIpvspQY7EjjkYp2fCPhsiVxGyYWpQJikNuAvYOCWGPZsyIwtWRhlpL
AzZZWmuPJED2EsWbJ552ngHIDlaHrWURrhInZSyheGvpW6vo9KLZy00zgmlLvXmanmTbTsGRO2Fq
d+lgPG1TrSmZ+43TqRQfzML4mfxSlfPguxpYQdxpQqFVODs8heE2U7BZKK3wQP+O8jk4HAJPq2qV
CTELqxd1ga+wI9ykIgbRaHBdxZYkrZQ1VNC32eGw5FCqyJC8E9sMxU5dmBcYUFPoHFjb+5T+AmJO
P5ywWbUe+NuJrQ5CGNCJTD4tV6XMfNmLL+s3TWRRhD1yNCxE/rrFOlgY2vjjC4CGk5JeyD/N2dXq
59xzeD6jIHKtB9a437iBbxWYjACmSyaqKnvdIZ+CsE+i56+me7g1EwUjSW5/tKzAu4BVBczmomMl
tBGOq+ZvHy8y8ioF+c4QFlfzMBFng0Sp5CKKoUgh3lVaDTwbqVfclD+PXq4GBnkdGG/NinLNFbun
AOu/7P3+Yjg1vGJsZ3q6g9EvBOvNVKifI2HpVS6GHB/ZG/cXm6tcqSPh9h3/9D05Vr2w0LMiEeOg
U4BOW8v3tdO3aU3s7HguXwSAL4Gkd7DE6E42phCSGavw5IP/glqSflSKE63A95aUtXowqOFi6gMy
ug6l0KtP5y44UqWZNiQZJOMdB1eGsZcuHuJbt2q4pLl6dDNyHo6LAm6lio0QWRWnWh8Kc2wT20dn
4x32nWhEBl+8i3xjc5APG87RJjzJFp760m7hSCCh5pCGDfGatjStq/KaFKD9JSjDBv1PlrPilnJl
ZJiVCFIxzxzCHcnvy5gnk/eYddMcJC+DWkqGfUs0h1v37iPNiKPrbP5cPMlZrODva7dwr0ct0pbR
SB1url1qElrHjhShWUcviBcMg9FsCojwu42ybBJBuf3XqgdKCMhApPwfKBKuDF7gr2wYrINKtHzF
SmcAImLEL10GF7a12nrM6xgGHCnvuXbo6x7Ly5keDlIrdR+NE2DWCmpJisrTYniJe8Ie2aQOGCw5
v5GiGVwN4Td0aYNE+ERvPVw/h/j7yMksw+pkf3L86TGS7gU7u+G+QQRjVM7igOQqLCC+ANZ5FrsV
XBxbSnMPttejQrr9drx2Evxfjol8hE+pBC0FOxpewIfnHPnmK0Qoyz6QeiceiCUuoO2gUq/VJZww
q1dKAvJsCqX9xWRis6amnD0JcOvn1P3KDIBK6LT8wpDDfgK/AIn7knU4nQkOxAJvfCMSzdQTobE7
Kc7dVOHPVzrjcg//gfs336+2bmYWG/+ospo7BKk8aOVZR6qeevdg7UERgPLE3h272L/VL8up0Fky
0K+H3xS0XXPovVMNCvOgnmnaX3hUq9AG90xNQ2hzAUIgASTRmkyn1W1EVexOAubibZI/ZPozhA18
9djpAegMuf9OZwTuyRB25Pa6DBT13xIQDWcIeKRnpcxy8hpxnXqlNSHDtBsyXE5MCCmtOf6X3KWD
Y4cBGc0lNcPKEWjbxv89/gOroy+ExtKAFfcgL4WRs3wvcSvjW0BRHwlY1LhHOB/TnZzyRRyaZHtg
/DeaJemfiyLoLlPNHYqjggP1UqgjbfiiApoKhpeTInuXWhWw5x1/T+YpWW/kGZhWeMdzrg3LtLSZ
lYdDYxTNZM1/UD/dULtLsXRnttIewPJtE4HKzMBfCjdPt9KQ5w0PdwvTXAc9bBgibAvOsYvaoUl7
vtQnN6qA1wPnY+/9d6V+zUp+xh/NKpz/4Em43IvtMjBCTZ6VdfIlA2m4vJFrHXZQesYvUx9W1A2F
fl0apBRpGZUeE3FXs42QQel365H4zTm+s4nmCXn02zPsdVvs/tDlk1CXf8YwIz0gAa8yOCGUKcUL
/THtQfJuoDtbhv6x2wkBD2QOoxe4fRDTwqOZBAbgG3qtqGPcJTL/KXccDNE4Gje/l8bBVWVvAfKu
UoBYabbplPsEFKrVOkG6AvXYRwpFJmxcd6p6mi8ZSrzEU4S/xlJ8dxJs9tEUwLYyvLS6jbfXDFjC
kKppX8Aj76oDwWUfDOgAJzA5X+sK/i2+/Yu7H2uiax+lsoRVlrkiglzB8etA0WgTaCnm0F0y20kB
t2Xr9Bk4YecjhZ33cKej7YeuixwBoD5Y+Uk2NOemGpYyX9RbC8AhmRlDayudEib6cBIpREYpJlv2
1wzpDtxQis/A1MqidKufVECSjO99WuJYj8qamydvsz1H2ZSX5wRXfv7lv3ieZfioFuMeZxj/HRHY
kPaHRn8tA010FDrq0TuaSPNW36esYBdxwbIE297xJKYN9I/ZlLxHLeir4wNDdcBKsEiFQ++jltoI
3AB+7XPlszGs8DS/xZQ73DBLyjpDa5QiDTjsWuhZV2Ltm3RjaOL9za13xvfYTJjx4GW0E9rpEnlM
2lBkGH3vSw4gPuPyWcTO23BbMoRmpyHhW95jv67zjliR6SkNb5z0j9SbAJTKtoU4JPr+I4+hZTEd
yEir1rZ8ZZKTFPhtnqpvVmIeS5tSWZSYSg7n468ZIzrVXGnQ/RfqiJCKtNs8Dsmp7lt+R31M3oj6
hCaA3MIPbvXsYwFeFoAlD/EBrj0Fb4M/sDQw+PK3JopmoFxP1xcbvd6DGgGgk9K/NNtINmZrmGpX
yFWDovTtVOoWoDPUVUaXQfFTnKyFXtSzroZr0C+aUq3SgQh0w4YioUWfAGiE/w30fQO2oayUCps3
JTY4JPHeZ41U4C7UWVf5AA6o36K1hv8I1Uuh87rSUDR08Q3p3LAvYgFYnx+RztJdHeEAC6hZvYy8
kN71atQbhTv1AG12i09n0f/EwCSTf0rEHsDYWeDDu4vfI3IzMdNjScpGIQBnByJSy8uj1eSlKjpn
xNwA7m19Bw2eF90tfWOcreYveqEnDb6Al3K4JgKpwUb9Nzg5MDektG6J3WIUwgsmCABixQsDJM13
sQO+VnX/25wzPWnMwMcAc2plKMU+R49cLtG5MHaRd4BVraHkK2HmMNKAQ/AJfNieJIwLxg0nILOs
RKsa5o3AZ4owuX0AXPB5aBVZZJcNvBfiInqfkhamDaoMixm/GxMyDEKRU93UVA47gRRYjuw4rKRD
V0Rl5eaqICgcDh0EJSOEyTlGkpMEVGEHR4t9LHcUJk/J7SzhcWY457JhwS1T2biu0mJSottZ0X7+
JLodaNM/89voOtX66+P23ZqGP2kii18vVP5F3VhzoKsPiOLpIme7wxtS5SY0m8A1l5OdRckT5tOF
xTVNl+gRcs2XgOLvp0Q/vz6MYA+hljJde6tJ/JXFUgnTDiosmBHhmq7GavVph23rCOMnpuHUbEGz
M9Ssb+fU8I3Hpn2Up2YMcYuPK44UO5F/N6T8qItDHSF7mfUabXRA557bfVu7mmnOTQzLddSu9zU+
y6dJ6TtOYgs27zgPBlj0+HJt1zwmdKYuAyFihOl8PzlNMf3nPhsu7HOl/YLYs/Y3hdW9yCjS/P8a
LgAgThx3jnvEzSjOg7bVrOicDWm+nSJV0lX6w1WOkkDnzhyVegoUfIRsuyGEFO4zuLhFE7OEErUI
BymHllqEL3nr1U3URH/7qSK3j6OPNRPbLWcdbiS0Ldha2nMfqLFjuEe7hut4kv3qzt3W433OhsZm
TTA3gk7RLBn5/Tq6Qi7XZK9/fGapt/hNPp9tdlFtXEB0ldQH9fgIYD185RyissRltrGglSuJNpxr
zX7mqtB7Ld9ixNWJzystyUcqS0ed3IQkNkCDeY1pxCVp4togDwhT5l+Y8VMU58/XkbsKA5mDz6yk
MdQ9T5MgQvS+ngrZ8ORiYPWQ4iqbzC3WAjooVpD41MG9vMuOdZgGX9D8ABnet2y86oaeA0kxHpPZ
lIWCXT7g8qAaAINREi0j/n7BLJYdLEKvhtcx9g8itKv2rBhtmTu2o1GFR3Iwb1YI0eHPsQ98qcN2
rElW3I519WHiA73nUMPSxAIZzuGiELxAmRlEE3hu3gcj9Le8oi2KIUkaOBTGkkCQQt07fLkUr9Y0
OWLato8XJtwN6ein1Iqqa+M1dCpMrIrGLB0yg+qqFKTJZzwbhhyMRcNvAW/2+mlExt+6EEXOG94U
ZoAbuxWyOgOahN/X4p/e9qLvNYTMbh3AjrXrXBFmknnlpVokXkgXFpKVUGOnixTB/dp3CEMwl65/
J2d8+5iv4p/10AjIQlHdIwvx61X34QqXe94E1+wcoeOp/VRCZunLE9vzvHAGS0Qd84MhYwU4R4ai
zx3CoqxUIn7CQqROIw/uR5YisPWXJBUndCLPyXCKJSfk51H23f1HUJDwEGzZibxqufbGwT80Kvhf
Z4kR11UnUaYUHNQAWNhJhXawnyzVYBz9mw/CWFI1deBamapSTFY09nEgWdA/YBOM07YgJRcBxwMz
rsvUcA0u6sIw3jWdQUzFyB42VYukY88hebfOCj9prIE4vm3HFtyagqNa+5mMbTmHmYncKnDyvcZE
wLxAeae6ZtaeZDSTEo6jzQOLVmT3DmdSDxsLscHeRvO2ANuYXnlvMMstf5/fglx7ReIO7+tsh5qi
wWm+XfmlD/9Q3IVeLqy3+T18tClVN7FM9wqdGbzIscCOMjIzhW3qsYK64JG0XgHpm9DQZwGebEB6
qdzzvQTpHU1ypLRQaHWrPiyrgkNsfjJix/IRTZ+pNqdmj158r61fyICtjq7IdwJrgOMbxCC4eyes
2U1RP7M44U+R1SSSwcE6YHMTVkv9dFetBzl1h1YvmG7WIdzE4BUOe+81+/XP72QmUP/T1uA1FLJf
52Sc5VvKjhdCqtDaTOXi/YIGy73MU85imyhLvgu2OA+H/h9aJUS4/ADCO9hQMQWsqXZfcEe2/Ry0
pRdpIUcj1RlEN3V+DJo74LGC1TLN7mh6mt+Rvg8b2CHWLiF9B4IJf5wGg3J3j1O9iTxyaO0E3jFn
oWsvIjdu8fhp9DSrLpiYi2k3Q/pLiRmfRPhP4nNWZNyYed7fMcSTSVW3M5tAZHdvVT0O7Q+DZbj/
9Misc8geCKynQlJMiVe9s8/qDxhwQVRhlzcCRLyUbET03MB9KAqrKvc27WkZriPzVTx1QVVcnKrB
wL5y24PMSAEdEkJ7MBvQP3hrN3cA1bmp9E874jQS6iRc1FDCpN2l9BFShL5sI6g8YZiors8fahXp
A6sj7zMn/LzT+OA0EAbU+weUhOz4bEy8eEIKIsOQMcuO2hz5hut3mN5umE1xyZv/9C7FAzlsq4tt
x7d95JZG3liP82bIU58gz4qSSCX2c8YcHwDsTVCOgY1pxuqWPlGxcbl2AsWHj9uk0uytsUkUD6RH
ipmTBNsz15VFOqzHnKmvnADTkkjhgSKGYJ6ElW7zZrtDmkYTfdeu0xFeHRKWsq7s4WKh+eS8o4R1
nLok8OEeHfD0o6KG97E/xevDPFKUlNr6timpJKYIhnfF1GVfXN8BIVXi3ZQjMhIMK9jFplMPrDJj
n5YHhRgOOejnTLsXmR5fv98wn+9wdNSS5EBLyY9SajJq79BMbo6ZZxiJK0qONCNJla4xh/EEIvho
Zr+XpLEgyKRw/au96vHnsVKpa+58jzHynnUreDLUxU7yLCmKxiLQ8+fZxL48AHdxNocIB/7lSzT3
mB0LgmsboZFXQVutFCFGLdMiOTJoRd+2s8glQFsPTCBS7x3SenfQ/9MOyDWauaMaA2mscQ6SI384
9K98TIH+7T55fIZPuPx59+cKanIGeUdnls+vMq6JYnqD/K7q2hejKCqXaHetWXLH4zR8QXFfybom
/BqnTrhNdhMBOsseWy9vcFqSA7itN1nGiO/vhuuDJ9b+p/1S/s4MTGZdEfIDNvFNqmnkLmCLI84/
x763MNFIviIKrIH06LIOk8zhCOZo2ytvZqsZzmyFcfH2jZhQGXurj6cSWP5xadd0KDC0sWMP+tuc
xkdMF8P1LxUFyXZHjhxKAuEej6QKeCZzDGKLQC53/sLL9JTPJeijpQlNqGl4qMwu9prlT/9pDbSa
cL5sno+7dk3PrAcLC3trLATzjV4BrlPIGp3p0w7m0avu4jTCrwJATmrlQkE72pGg7QplNLDg6cub
oMkjXWPqcAzvy8X1BbNEZStGsLZvmtZhla1zhBuFpDJGD/Qd7y1kSaHYnBcxFbf/fT5q/r7mNvBO
OkeArsgrMC7L4JpgcHnapV6439K0brTA6hcjg0wpEfCc6hw5bGaBZAYq0zC6oqUGwfCfaq1HAoGx
X48gbKoyq9HYDV8W57YjnF7WAOD+uSLrW6vEEIuGrgkJn+wdcaDRFON3h/QT0TGvYBnZ1G7qMVfk
qbpzgTmK25XesAFQRPD+yik6qmuLLrlSGcmMyKyrCQY3sUZpHal6nwcUzP6eR3J9BFySD6tpZuTE
CXWq5ZGirc7yGSXHGnLSOzYLeWWaRvriCVmHAmtzUJSl5NLlooX++CzyzCWgtcbwLidEo+I8iok7
xi6aVskbWFEqY4M9/zVfnZCGorVdvjWccxUfAoMycO1WS4TBWMrh4G/bpCSySQdusa3km8CrXU0Y
9RPM3CWCYOxG+yhlDI5c4K1epmJeEPbRn3TozvFLQHaCq674FCezkJ3QGiWgYUoucmTBRAPz/6Tb
PzmBjJr9ZalEFJyvXjxn8jnNxdI8bSNyCO6OZsKgbQFm2yaUyRglgxuyjletAkCIqinXmT2b2ld4
5iiaU6UAYbH3fSVc45UPans+YBDLKQtnmR+OX7qtpxKyucKaYatDua5HnWztjwWYXQMbNl5YP5QU
w+AoH/Yhsd+U77mYBywT4ZTxYeOOHP1h9yw77OJR0lk9HaUe/kTc6p6PKaXRVaohPcOpX7niZ9+5
VVr/fD7BZMR/2cw0ydZ+kQx8lyaWUP5liptE86tYu7k62sg5p2pdWz9ZqdPHRQKG7qySbH536uou
iXnl1lEwqBjP9tZ81WLsT0zh+nBFGIZcVuhhP5pfkGOBFRRDzM2Sxj9NQQdh5qItaaPQkOK4gSn9
eyqLxrFlkGaytcouPXarGbyEWkPM6JrtmpimeM3HjDntrlaOGlRhDDi0PXVxP/3OiPZaK0NqXfr/
fVQaPBkP1JoKL9xPv0YPorwzZR7onz1lA9lBrVvpVb9LCHpVmZF6xAIcf1Zvb5rJF9efPtivcUqO
EKjJGdJC9LieXMU+yhquqHqNuateu6gWFoF0slE+5uJmheiKdqfb9Sq+OgBym9t3M25Dqlp4tBrx
hnDDifwCiDI2yuJm3Zyy2ND/pZs6g956UoOInrF5ijCUxLX+RbaHzC/k/q/ybwj9CXWBdnBo7Fhc
O2T2nmRRJJJXPmrIKn9OHN2gyzLr2/q72TNnjwn+BQo2o5XzwgpaOqGFWEyEuV6k9jtjH0eg4Fhv
zqVfphi+89yK/FBVk9kjja67AqNUqYjDoz0DCoJdfmWmvfN20IZkZHL4hNcull1zIptkACjKaTcI
FSyXZWTfBOM04hAW9hDSKq3zZ4XuNi/O7foUHYX/OH3KU8hHzy4by6jYyoNasQhGgRWuoUPnZb0W
5SmnuSBCTkqWrv/rnBsb+ag23RrWOKyNaEEU/6OrV7mjo9K7kNNPS2BQExV2bJxkHL2pfe03MXky
IisaQ2X6qLsoKk7zp7iLjFoPxq3ri4WIsq6d/RyY1D9EbWf2yvsGl/fgFtnKtudT/UWKFwjBQxsK
BeJNRKEiRXMxxJEop3Q3fIX6cHCO8ddM2l8YWfP7m+t/1g/KHBMeTDxVQW/czXgOAflX6cgIJbb7
02xA6iVQzXGFxolavdxWVVRFr3f8w5M9Q1gewUum2zwDztzRzbZAOQqfkZdGAm3zFIekT5aisEyp
X3ap21WO51hfGVYEACqykGxLzivH6mxDk0+orOQc0OrWtjs+zQMB7LZeo4/IEo7CNneKTm6JOuyn
bw/s8eTsEAlAAGla7BtOCALUZ1f2M67JkNZAZev/SD9AXrPfA7q+/kAB6Z/hXvKbUC9JMvbKY+nF
zC9n1vi/1MxbyY9upAEc/1XYulRwNn1b8DmxRXSWOC0qo6MpTjCFOLUR7REd/6mKpMhqCvjr4bkf
685bFvGA9WZ+J9Lbb3Us4TefqVqoCiZUPOAACj3e3r8GqbsFXI+GvHDSKauZEtzzJFv0riow6usb
L/lV8E0IdczSr0bND2vUTbhs95zG7VJ3yFPwp9izhJcuHz30aREDSewsWeE7cII8dNl7ZFwPQ+nj
MX7BE9kMbMHX9qmKt751cjESi1REnZLRB26tNdaEX8EkkrrMIHdmAFVHKT0MMdYYGuzAC7HxACMp
KRhxxxhbeWOaZ1DQB9wgqEU8E9f/c0/yPzm1GiWDju1SHQSQdMCCsgKEfoYmRLtEThusEaDFW1nK
B4AW0R6nq+iEbgqd09oNVed+2xLqZuAOjdiv2Iq2mjA8cp27spn85JLgLdPNH8JSLluUv15StHJt
Uq4or75BAK5mhln41R5sPOkynECVl6YyIYR0cHjqYN57XooHUhIGDZSY/VGoOpnbXVlG6Weh1LNQ
yc/qxL3pVHYpkakgk+72E1sJSHTipCrClpfC+GYriGXjO6Nzyxhhu7U2f9LSpobVbmixS3+a9WWQ
oB3Ea+SunqxxzS2zdfmz3JeiQj7vcGebt4jTF6vAkpBmqaotfLOuVgQZ2sIfv03p5xdn5foCsBCa
xVz02lV+1k9ySmR/A4QQ3OmZnqHg8Wmy68uqOvuXAAJmX2XtxieGJgW+g0j6p7kkMuwOd+lqNv4G
xXIGqmhTQlJ8A10W7L+UzDjp0jYKQOTVSWrEH/bSo7gZI0UgWX3rZa1+z3p0mUO5utRYPjLJ+E9k
MbnLSWtl9pvkR0aWpPicNDqH/0WNqNp8/PmJ94mreB6kJJmo+GglJXFcwhgRgbEXiSxJeKchqWZA
AwQdqPutR+4UD1A23DPLPMRRh1YRtUlTLPNRUX3JzOs9o4kMvvmYAOxf8QXidcixrET2CIj8tw3s
MV85VWQdInHK76K7aUNLaRr+8UGac2uRM3jPRrAONC2u3FJgqKlyWi71PKHuDkqcuN0ExSLCB4Po
IlG96Ni8Z0gDNEQ3YXOdcG10cv5uwjC9BT3go15zlkRfuzWYFORqLYZu+G0y3wSW5oNJnot/DhsS
3iKWFD7cGhATLgzcyhL8uWiREBHCdpbvq9yGXMZHHx2HyEg3lsI2K3b3yWabyoNHoOJMO/96ZPl+
WYwgnGbY1cxi6pXackOOQUvaKKrqXKHZwygQzTTfE5r+YuoM/A3zVuA1BfNsP6Fz7kDcPv5vVG0K
VjcHS/tY8JqF4ZfDTUkE8yTC2VVqxcj2C56uFYg0sZ3YICgzmewJrRmGNCPyJlupvCkymNHcrwxB
hyfZoKmkagXomrXskb+VK/ptZh/T1uBQbW4qAl/UJk+JbAjrcgJai8GH+oepOrrVd4TpiTkX6sfG
u9UgIcuWlwNbndIaRVN55aiREPNjkCf6zXy4ytQA+Rzv0bftjR+XskBcfDZpn9Cv5oI3SncBeja3
nX0ou85lQ/JiqeW82F3s0I5cwXySMYikDmW36SIfPNxzLLkDDSEUmqCL8jSQzK8j67UfThBgaAY7
fsDlP4GHa6gmhk238vsenidNIsLMYYWijMCWvKgN8N7i/xJ/m944l52RrcX3Vd6qR4otL3RUYGnl
/FVVJngxRtT7K9aMcfblP73z1uIpbWLK2wZJ2Q8A9IPJjkeKmOB5awMMLkDyLUZ3lzp5UQ2jFCnD
gQjQ6aEDBti2N18hLjKAVCQ2HMcY3LUh6Du5yv/Lnsg+IiLOh6lmAGcxnANC9u8/TQNLS8AX0xOg
5Eni5o6U+BowJDXxBnxJMgKuDgf1V9VXqWjNEnMr29fNK+zR1j9eAKaT2ZlZMAc/r+svecj78asR
he39WdTDBwSSeW/fCKhiINBiTT4GdMcrhSscZjBovU96Bb51UBJRfxIIfiSzG4/YjzyhewcmgiVR
ztJbJYfa+rbCPTNYQmAaayK6mlOS1mlwk43j/XvKIDiwBRMa9QODlPaXzVkEEDpDyM6IQM3saaxY
q/AIfd/MrYOIVzyXmx8EYaXIIf6gxFQFD2Nin96HwrtA359YaxrWOwmcIiINhNlqYov4mKC4jD3k
wMyyFiycTqxOtfOJHvnf0MQZqXTtku/57EzebLgaUUAIGz1HvlEiH+w0WUPOVe4BwZXTe0HDzC3v
B7uQJLa4EpANOD6LMvfgLiZzq949ffBGRFx0MUtoKFZRAeaeVO8w0tCYW/HolRxtzpnuR/O3n5Se
j/oiAMJz87gz7GtG1o2YZ9Ik1AUSKM1G73iuCqo0GxgOpIDWf5P2F5C3ZovIF90g6xVUIDuuzQE8
jiiUxH2ikbkkp1zOaU0Hlo50pEx41LnSb7FdJW13IDeh8D1e1FyqzgTa+iuuKTdJm/2MTZHI11RB
L1UKDWFHD+f2fnXjQ1pNyk16TYIuMTiLB1/TtM+RpzMkRYuDZ6yETjuWAZlh2B/vfZQD2ByO4Uf6
FPs3lWfz/kNrhZj8cCQUSyEBWxYRgCuncskRqpdyFL7yVfW5zC+FTQn3qJt9YkZdWtEUou2k2koA
l3bUdif4QvNptrN3z6gBQrq0dQR58TKy3o/J6gsfnqaOH/LbWaoSoy5w0HsQPt1DY7065rtcoMqH
svWpJsKKcdp0mrwctUGqJCfq9WXdoZ+H7Ddn2+V4Be9njSAgVzmqwEh/EKduVZQAZON8Y6qLQGHM
EnIT4SIpdww+cI/Rn/3FNQyIC5TsZw3G2fls0fsCsDMwstsc4Hjbs8YzsLklKM47tR3XaZSeSvsO
Dc3du7kAoTvPjKFQ+j86FAlcWK7gcX4ME/4nrXNJSZD8umaRRq2S/2qleaKsE6wsdfqE0zAY07Op
FAIx3eNCJelXo2gxP8qgkLK/wGj4bJkaMQxi0gbkcdDsWKY7KIiUXlCIeWFFWlFRf2sCpynZTvJC
j296MGQEQTn8TbO5YxugkRGaIoCAXnOp0XZE5H0KP+YAURTfUGcpdUEXhJlp3XKLL8oQlpgEo+z7
jtNYCm9BKYL0hk1I1MuBVVIBGZBUD7vy4EZicsGODRWvbCFWhB8SI8OOCos1EqskLhH1u7+QWO4l
2azTDEXPLnpEw9EeDjkjuvN1xEHRjEDoiO2qCA8/g6klpDlgf7lkykSwiwI7cnkdiQhMQEFFVihs
dH1r4wn2EyXmHiKFHSARcxlzSQ7D8nIBMa5zvPXJ0BWamd823GrkYD11PxMMLKQzab1z33RHgYUt
xvDkzo8VGfN6xBcRFc+D6uBiWtPdg7OxLDS5LWzd8IGTYp8OqSqGqV6pRi5/3Szq+B6RiDazVltN
IrDE6TekiDrsQumVZXlFMwu6wVzyCpzwqYYi/89BKe/Nt5y3Wb98oqZLhe9mcvCGlPl5hV0L45oo
MhqQ6YhnWPtBQFptrjwcNs4oz4Ns4Ed8spqamBOR3kdbcR47ejZDTUwkRDkltmc5GHHBqudwlWyq
2GF2VYMBL7YkQaigB4cRhmQK3Czy5z6c04srhi6ydgodEVahSyMFbwmk+QzOq0YAuQzf3dcKQA5S
LBv9maO8orkZRFeyt3TUbLbua/n2qeF+IHv6lgc2TTyZVEg0avFUKf78+/Ncyrin/3ORuuMiomsn
44cuaN3Uikip6LbMj1IqMLGRY4i9P4xlg0IOD3+DXTjUJeKlIMoRlpK+WSZM20nmCPGwhmcnn8XB
vOjUU5HzJ/LHw3TFb0unhEDiy95hQYFvz9sAJPFGncn5LlRKPfSmxM6l674E48MMLcXqEvkspaOb
Wcs0dLUOt2+UY9JrnSAn+l6jvF0p53FteB4kyp5f7ibZOw5dnKsttUmMJkmaTwpmoDwghJXHSCY8
YtQrgpCjnhL5KdlxoNaeePvdjsPlABdqrt4iQrSUIqD2MEc9vWNABnwMryMq05m3eLKkWH982eOs
7/8Yq56rsgYiDA1gN1s78j8zxmubMf5/6n28t+weiLHi4c82RzUw3egmlVRbsrFjqIy5fPxLaykx
T21ixRz0WpnsSOgh6v9GiHcPOMNlvcb6lJKCOZ7zE3TQZImQkQmdYw1wXJYW9QphJqq+nNime52x
Hvk16VQqo37xzp03mCgvgptDrq6vkwJmk4DkMLVUW47jBrUaiIGpVh+6YNVQPtf4/j/O1U2En11u
rVyvpr0TazhnqbQ9esSzUFzC4qm2Uvpm+EPeJmECaK95PWHy/Spec/Pc7Nhdtg79DctjmSB0YUjl
tpPnPRRZNMGsZ5LLhmZLc+8TrmniSFHrnkrThFTFZ+5Vo2HcamSNv8MXPDiy9NUTnSxYhXzRb//C
AqRv9oPZgBRp3B/gDwBhBJEoL0rQgJcClFROMjmYSg7uvnUH+qsxBlmo1oHZ6viGs20V04ZGzING
J0IxTrkIzy5gEDvWOHmaBc1S4EPtnnMy9I6MInoec/D0F7nwfGTZa/fDZDY0qlpZK+c4QsSpcdRa
wN587SfrnRjtmLCQSvjB7/V4/B9/dWMXDVdGp+/y9ksvN5TPZYTh8FEPYw7yjEzll6MLMAx8mYDU
z0qQ9mXDLwWw8aO//k93DkY0G6Z0S9TXQ2UoN3nWOvQXg3+1d1wOYDiFfcKFULiy+cm17XHyERf4
v6MiCjHH+LVPjNOI+Y56/JTdIexqdgBRsVPpuq2pVJ/PVAw+q+4yQ3ue7yPFpAAfN7w0qrMv5NXQ
q4xxbuqUXp0RiFP/rdI0RRJxWMsfKoWaBuIgcw8MvXLHh4PPLs5sS21b14R76LAUvf+9VYTa1fyA
h/nebeQpQVF0g3i7+Up6UGMdGYBpBkJPfaHH99qPZcDK2OqUOAfMy5LWjw+4SFw+2jeFMyc6l4WW
tKEPErAVsMCnGgEyvyetlTYeq7SXxc5pIv8jTElMK/ndhM9AmmvMR/4CAa3FIv0caFgGV36A5oRR
TjZ5kyILHgGFrTh2JDP1/aNC44Yc8sAbXIrp5Kc3uaf/0IOcrF9rt4DdQiKV+TqRJcmt7OFVFe8F
1mjY4bKlPQED6HUWtCcK3yZXWZ4YbiHEN3bg/OScxrA32f67KDrbkocZohjTwqu9NZZ19SLF0u1I
WQDu6VM78trXoSpu43sEvJ6m8J7jNr6XKtQuXJYYbGc/MAMsuWZ/SddkKk6wvMQ2w1P4KF/SdzQh
U3dZ7JBLvcNtPC7U4FOcNhIMLqc6UoTbFeJrj70K+Dwv60hZc19BzhJTnOyolkmYo97rv3RD/w1p
mYiueP3CR0hGz7njFCMAIoRst+qnBf94T896jMOootpka5n4/zX0LNVeiU4TbhM2Qron/tPQvp7D
JaFPBazzciBBq71QmWLgYct2UciHkz+YskWon06TJkw7AHifwDPFTbdX3No+bxd1Kd5l07UHI9c4
iwFGqyw16dPng52n7S2gHjpI/QtNzOi/B9XI+Ic5PNx/r3n00Ma8sh3xWCur0D5ivT0EUaJNt1xu
OwEaRLY8/2I3Toux/AoOfrTU0iiJBrYfN8sjY3oRQ5EeWBWE+qkEF8rTKrB27Ha5eOgltMkTyolk
iwkOhDnHg61NNCZxdZfd0zgvaTNAtlfPRlF5q8Zi4bGNHL+gaX8Ba+t1pImgHXg9z2yn+U2WAga9
HOj16MYGTEIgqPanyGc6+YsT74cCUZ9DJRGF0VDLzgeofSVNbB8tpUHCo8a0+OBCtfYMlzxqqpx7
N50Veohl9Wv0Hr8pzE7vVCf/MNGTjST8z381gObDGa2iLCUYmFqxZkB66RrnFbKnHDcTV242DPAO
X9Js5IeCFQtpQqt6F85ExuRx8Ee3ODnpt6GDX9+5FIR9hpF2AvLG7TbCW1Y2pwdWuRVL26IdYCkL
J/PU97W3j9WvtkVNB4bZmoyYT3Attq1KohtiiDrmOEnF8JrgXgwjU5edOS8k4MIlYy7cYkeKVHoJ
dZKCQ45L3ELCplmdr0WrxkTsncHUjyqDYbV3mnBCPpaNyag+smERMY0rVe+MWB7dTa67LZwjxYXe
t0h1LnQZpWPGhM7TKo1zfccCGTVPgX7TD/tp2hLvoAY54vBqWWnb3OJHSlbgQPEQJyxxgjpi1xbb
AWLASZegDp6juzLwCivZlN0Jw5h93P0Sxz1mRspFcMHioDOWQx/Dp9KEa53SJtReiY9zU6VdNFYL
SoAergl9GE+8BvyjI24yja/ueOhPsX8CVZtlXyE+zct+nEziDAVmWkCFb0SJ96T4puVpcdYakDX4
vywdBq38b2B003VeLTFuexVwq7rXzEeMrs48A6WA+8vOOrn32vf3Y5sqBVNJx/ZFdNg75jdDcrR4
12Jhp2TXugqG2NvXYTGF0I9uIBMTGtzfxzDZi/5P1iVr2GrwSFyUyH0Jl7ZNIyfWxosncPxP3Q3e
YQ+Y6J12dNmCTTi+3OJOClrSGxABZlI0o32vIlef2RGwS7QY5LcGBnx4d5DQR03D1x1qXvrbyoMX
/Usnh9aKt3BDWQ6tkHvIJQwRtVxz0DvLvXUnNinkVeVb8Pm5YHUTtvD9iFGeP7PeVTHmyjnC2OdU
1k7cPYQk7O1ZLLSgROvQiaVTUe8eBo08bpYhXaCbyffoenlrJ6zeoGu5RPkb4DaBIpuZi7/U0I83
kNKzTOLM+Oa/VLh3i3+p3/dzbQjuyz75+LA9NGj+PhxcW97GsETIWXb8nU7JybxbTfAmdhvzsScw
8GzKCC9TJ/9qOLpE5BuXbxPKJqfg+FWhpU5I6B+8OxyQEbHAZIESBk/lhmsM5sBXTYTM9duEYanY
En+nPBAO4G7lMhS/XuBPMj95l3FpdzU2AbQHGL4R6UOPGRs+UDEOLLm1NE1+pNoWkKUnWVzm8D/p
0Zf6tnxSKBntrnhNGcsX1kwycKQksgT9jZueFglmYOZzrf/8jTAr+ae76v9dsw68Ttecfv4FPUk4
4DLM2eH6p+SAFQ8wvcZuIRIMDM7pdSalYqe/Bs0tX1RvRjmccMMjAp43mIE295Ew9w+COcW7Mjrz
dYCwiR9mJq2JA2Adq6NL9bfNR3WoUQoGAjHETHjWwWl4j3kPsrypSFfX5+2SOwLL8WDESvyEFATF
lZjwdWaUg8RlhnJQlGREnIH5sZv+M6BrC0QVzVqkWdVSiPXBU3uWjhCsSd3QPKUDqh0W0uNeJBfJ
7urc710nM0WPG6NKX+KuqesgrrknqG0l11YnFfct4bdb3gueNlI8Yfo666McQnX2Huc9vRMhsePY
gWtQbTel1o6YcRZYqe1TB4/aMuv7o6SUcgrzJBnlOg3opcGbE/k6UyJzpH98IuhtyWcfMKJBArO5
zgb/5oj7H/KVbOy4i1THhtee9PDkRGj2HCO48I8Q4xY7uT+oFoj+Fh76Lwzxrf8PHQ/2W4VBqlbB
mCjykGLpxcqliCgEIitPm9Z6aXMEB/A2Jhnc1F64TtLzW2dd3NK1uFL5LF6rn7cFl4eNnVfdSHBh
Yp/PG8OafQ0GhnVl7U7/kpMdqqGrGd/MAqpJUbRsX19D+yzxRpwAFTm0UqhbuLQt10w5+ADljhRK
2BNNW64IPGy7cFkFEUtTga/dpO554zdcJqiFsQK9nnW/EYK1D2pQC9vJGG81R9U1a85cTjBG1dAs
ENKK48YxcZndkTd64QnSmYo107RkrJ+kbJaO9Wn3sUI0lC61zTR05+nW+/Mp2qBfsV075LrcDVk6
9Wy3bn6PFiGkQsVS+hu3iVdXd8Ld0jroxjmzo3nBoiwwhPFPitlkf7MlmJVXUWXd/3gIsIc8RS3l
dxHI7gM4s7g1XpDUFEpJwWAitPSomIgUq/k6Aso7DjaeUUuOOnWqqPxUS7+7Pw8yQgNV/OJoue8w
VfaDqc+XscuKvGRpr4jqKixUtGm9wyVTejt3/qV56bCZzaztedxj4bSmvXuVynjKYrTCVD7oyONX
xX0DsjmbSIhGCoePIx6OaPxs898HLRRR2oWjHN2Br8K9lLAhBu1KatrtAzw7RUkmkVZ2JQgqDf9a
W6pMWhcdj2rLDi4ePQ/uRx56YScvHTwIndncQIr0cSg5pI+kI0X0FoXM+iq3Trnkuq82kmOSb5bJ
mgAX811/k2LAXhdit0tfF9DbWPhZdt7+cfMfI32wqiA/0qbFmRBfyecFy3GCqFppThjyYQKnihAS
CYMQ9rGsQaLH+pO/WJBOTGGb9kXNE2l+ZIu3dkGYOuev89kP6NroYHH6x4NUe+urE+fbL5frrzSo
feLXX6SiHWu6lVEg4IVHI6goJrAmn4vKP12f8Img9kzQMazmIhVvJLXKyCjFk9pxhIJ6y/jKUegj
D0Lo3OsjWKGMVAdTYpkO1g0pV4U1KeXYWo29V2hW/4OmSpw9o5hwo/J0pUkZP/kGlmnftJkEolcS
m87zpuYpC/X8266Q9N6pjknXZZrHwjxshvhIgC3u9HBRI3GUDKXo/8UGTpgDPDEsxaFBn/rNpBmB
niReoOq7Hu9ZmwhbaXaZJtG5zcRQURlsfN0U/9aOY78D8k1yAl2YDCSswVQLSH61mDkBqYn/6/Nf
jkVmuXNEPh/dCkAB5SnzX7twLKefBgUf87c6XypJ6hpzmFknM5fysRuPwKOMj8ulNnVngd30YWqR
Zru2A1elSX7K+HeG4vGMBBudYsgIuEOoB3S/TNzf+zCCdgLOuhzMzSyFfGhdEFWfm88/xyY6/H3u
f9ZpgQSa6RZNk03VAcoeIQKCCrV2KSBTVqbpXhqnZY5VOgicpfhE2VmR69/Vc00iUQaszesbvawt
BPT8OlpGy+Hb48C3xGh2AkcEiPkFZ4HE+ySIM39xeTWEhSfvzW/TVXZsr0tESWFlksx5NVWs1wWT
mAXMjTqgboGy3IjmE/SYWJDHMBgG03y5liAwv5Q9Uz9AjTp7dgBmdIjAUCLlB5qcJlnjJf1Z/jWA
k5mtsHwOz0/shAwowt65BB/46lb8ZuDRVV5Cod9srnIkn5Zy+voE6BM61kx96E/Yo1+5Nyd7F41w
tgR386HzG9gkiKUCnkJuPHQzJSFhRwTjyiQLrFhC7ATAdWyC6Zznz674WzE8aqEIbB9suE5ONK22
G+yEHCrYqPVFKrOVtkWTNWpmzr1Da6xsJIkTpcrr1LShwHhQZamYUvSh2CtPGBC9AZAbB68LJo5U
dXy3UFX7NfHdxRTEH5a1CVyyTeyXlHIYtOH9nfZ5lTWahF4RqXfaSd/ZXjQ86CWPE78+o1n+bx2+
yNiinzvh7JEW25AEObQn7lokyjeAc4nx2Rhj2bPM2Q3nzgH8uaCllVX6Z4pOS8rrHwUaYINqGxxU
pQNNHgSf5scEMHWI8cC0yg2YfxowWhC5CCIvAQCCpywzQdCAcHePyKksUMezUlMis1drRb6brgAB
TPzdtz1e/9RuRPNlmlWgs1bqpe9xWu0omsuCaYIs8Jo+avmBPAxR5cGxtL/R32e2FE/b4iyRCjFY
vJb0uMI87NVmbpBTLm1JneylxXnUKpPfxKx9J1jGM2XefT/CgqRYlNozeXoMM5TKt4p1u6oAwu/w
HCPGbmwzevF/3RT6VtV8A9V9hrUk97dMGbMEcBgWzJR/GDMGYkQmsdTjJHmD6q4v9MIpjlO+sGx4
0HknFb+7jTKNEcIC83OKeUK1GistsSyQUYjzAauKr0H/U67GJgngR5KR7OrfnKUstTc6SKnFBwOi
ub8IG5g6G9sAIAFdAqYpsdSQyhNo31L3PHQniYdHkP8yF6Wb/sfsOXz21ifE9kzlV7Vt6XfYDNCB
4n6JomIQs5j+Pmc+7OLtmwsSv3CQx86sByvO2N4LQf9gj4Acn7AdjVY4Z+Ht6RC9/j8lQoUy8Ugs
XHGhTKEL/04/eZcgNHjxkLpwkpkON9yDw44T5BMhPNWb+C8cdbvXZn+ktTuZA3E52aG9E3U7dvq4
1D4r900oObzja1WkLaNTMGw3jw5GEZhpaWL298voQ3y9PZccjZrj15PGqXs+87vNBZz1WSmCeyMG
AxreEyRHwdPHB7lcAgxyH2/00Yt3vjZPqQ2HvAV/pyIhd5XMy8df024VSVQYM0DsfofGkT02+F/9
sAzIwlcsgwSP4t64Ew2XfTIPuhh51ah9tfc42a6uXwJGHnodsn6OXkms3c+CXM2JjxaR1QMo9kjy
i+6nOW5H7EzSeUpBY0A1ID1xNDxcaRzaPNUHCwKFOnFJl+RlPN1XtIXBhSvfNJ7VDIiezDOFELJC
iqrrMgNQCvIUJNJ+U05regqzQgUMy/8aufM9MqkNIChoSZpmokDmh14h2ubi1QNAG8jrnPM1Nf6n
dtx/GHP1iOhUu8hp6w3QVTYyGXM4ebmsHCKXqC8EAO1UJP5G0WpabmHN1TTmEGyCFe6gZsmW6rFS
8Rp2CdmhVblSA0fhzFAwuxyGnXGPwOHhEzN/UqWztURrDb+aWO80sbEEx50IzSGDXcSqQBDQfVE+
wUJdnW98GE0HUZDEcqsDCHKrIu6QnNCLnljzKvB2XYy/FUBr3NxkKwJ9tVINBmhDjT+3nNHfEoXR
/OJCnFIYk8A3LAzHOpSkF2QI6P1QoRHT6jv4QTjbrisg1ZIVNYvcAlEwl3krbKNVH63ukaEnN0k+
d3brYhJuEbFZAqFCAxK5XqHinaifHNLrnjN+TJEtdPfeIEtcIy84lD9P9FRCzIEMM/6HZoGGU+dO
j53ZWqzw9KC3FKlMHXICL8p/QHDp5d9PCNZPn/N2MEVVT1tgskRmuxps4nfTge+1/93/Vc6qswqT
rsZItMUD6ESMLQtylOAOgzzWa7CVbGOfVQngKzcctCUhpVebjF/46EfNyeNqRy3+/ocpbWwHpy/J
fBFHdr/o1o1o2TXfAmTNfR2OxfEJE9PtjY9ro7MYJXwqBn4/+efkX7Ecj43BV2cPHgeMorPjyr0b
RvZHt6SPtrHGMI/pciVGWFSBGtOJkfhf2HqqbGcJi2f53VvamqUaSDyo072wrYJSo34hyM9c/zN5
A42jYnWa3t/SJ763Y/nEnhGpMHzC94/2cJzETtYgPuonrMcEMFnIGguthCjQ+wrKFfGqr/i1dGVq
71dQpckgco0HB1Lv3hZryjO1RJKuJc18ZWLlIoBoyVTRdu8PmdjQmleg8djVX7PxqOpnn3wNK7sT
7KFQ7zeBE6uLkZSXrKLWQfQokonOMbvoUHgLgH8FLtqZCYkMx6ulf0G6fS8hLCo1yWaZ4j5Zv7wz
lNSdp0m/PcZnL8+Ulo+26cn2dfl56M+rmiRZG9thAbzz2sUQpsD+pv+FKk6YmfKM9d5KU3oSfml0
64yuunUeRpkFBL2ijbBaZRCPmh5w3j1dtLhx+ju7FBeaSwcmSgXHAEwsfR1T1FDzPUbNpSxhONh/
gT0Vx9dT21IgCvsIgXp+4JJKHHJTKfiSzm+oReGA1UhvwyIKbXE2hDXTtwvJqxN9TOTmEQCDSGgu
mn29FJsL9wDhjueiIs4kgzUTgJY9AVnK3rD+FY6K1XuAmmRBPRBGrX4FWbs/thd76Ls5zuYUhPMw
90TRcam8umkMa3YoLHv89n5VNdhHjcPwRvf2tXZ7h3zJZ1WBQas4522n2Oq8I7Y3K87rVksoEM5x
MC3YPWv3rVMO3covb43VK1V7OI7qJ3bWrsZsuCHtEySQFEDdEpaITNCTdyZNDj2m2VeDpTUbpdHD
pmBWpDcp+3Nt7yOOtEeC18Rx2lZgCdTmPer7O0HGIFdNRyFCwyVDIUXkrs2/JGqB0+utG/ZMoqmN
wzz0D/VNRNu956c3vRx+T9lHtIBasnJuXrf7kuATSlzf9Q9hjpMJ8vby2d3JfCGNYOfD2ry7QAnV
HL45aCg+JE6N0fYtg1xVsOZIgeo0U30byFDjIiEgOXfFjc00tIMr3VzNPaKLuhnm1KYvyJl7/kjM
NmHPd44yX2iL5DmfmKSH2KIMM1iRCzXlIp7plSkb94vrcZWMVBJglhvOg61dtgpThMCogmCIzm94
DG5YI5H4opJB16ktN/hK0Q1XQKGBfnS2SSMHlu0uXviec5Tv3nVxGaNiE98YLnokoZnHvfl1uqbA
OV5zUCKOniZYCdu4bbrRuln46IOXkMUNhd+4UKpZ+sqwhoi+h8dlIAjtrChHCBLEbCjEBSBaUG+e
JBmKaWqhuZ5LYQ67LqqY/zAmmbsg3s/OJldY2nALjnSoqzxjtlCvZZoucSNpNqmd5k1WnV4P9RZH
hzMxqJiG/7MkU6JKk/qYE47Gr/MM4E8S4ujSUeSPmBptaXfEKP+ybLHgEzUUmYlqigjjPIck2gMu
2BsTcyJ+MJQbo3rRHDfPs/qPmucwVi1IMQM01soeK+nDVqofovktn6S0d2GH+IzNfJWkzIscrO8W
V2pdhL3l2M8YExwxprkOQ43cGujENvmnhbdQh7nOnCOmjv3TywbRmszn9pIN9h1q+xWVeQM+7aVZ
+y+SFfVlp0SbEeoCcb73ua3VN7uR3LP1Sx/ebQn+6j3514733VMIB6+lohcmBw3Kv8OM73dPTy2E
i+tYCj0FpGQLG4TDFqoLSNuD/h0EBbuC8ZKDaSaRxTfGR+UGhPLLbrReuZNah0WFSpAEa3gfNYPH
u6LiaZ8Mw6SHoCpOSonilkcCOf30NUpX7ltD2bcrjyZxp+Hyh7Gm8t88psItnKakaSdSFSHU2+16
+CaIQ7FKLS0yBY/VdXmQm+Lwt0BCG7mGf+oRQfrnNd0nWoFllZcH77vinBsCWzL2gAYw3W1Jwsf0
VKPj2dZBh/PUnS/TXkwfo6vWfqz1RnmuT+phKJljIPioKFc8T4wHhJXhQKhQnWUITRs0BmtZTEVF
mKkNrqrOy+BPrjmfsZ9lVtVuFnhbPIO4lJF3aIMZTdnySWNRV2wHCD5hJBxG5eqXtKNgsQjmNSnv
1Uql+EX9xvpQPR5C+vk7gTECnsHI29cAPdFXJHW3Bkd01ERI2TT+9kMb1JxjOizDbmuyd9xabmfr
+c+WcvJRp6rZDclL+x/IdHlgbCx6KRJg7JIbARgohbRSLOrCe5kjrZvgC66hcLWBSBt83cpzpD57
zc9nIkiIYnIaZ80vXilBBYNGBWvTuzgcy9WUbmUn3A8dn4ZnDZ2jjZsbBY4LQ+4zIaLKAUXAAal4
sHhaS1hLd1C/0TOCo8ijhbEo1qTXD+ar2nF979bCAdMWmFBNozT0T0pSm2eKno6xgJdJs4xR270c
R2G57jA/y2y0CFfpdWm5AzXCMQL0DaZtRaTiM9TKuf98Pl5K3LZtmDNMhf2Ubmvhi294ohEWbrCw
tuLbTHdeFX4bA+fe0X8DKvZ9KUjmhdGR9a/ANtRE9QsH17iiik2nHXIHWICIDzy/kvYidJdlHVMo
h9+9w0xU/Sc1+AvlMmBOBt/QhRdT2MLyTKFVrgs7zEZ1QIAjwC37moqPxLOON77hLZ8elOHQpa+C
gwp0SFIAPIX2fDMMnJkYGeqczIA0gFUu+s+If9pID25nn6/gRdsuh5OOmNi+jHzYBCzpHTSIdq/2
+QeUyb0dOnWahTi210SzchBavgs9ddHJ+iDso2rssMe1KcTj9Z/bk9LTf8+09nV8kqEYnZe2e33y
aJ4VC7eL0tQTFlbazduUqUVQhbLQevohPvk5bk+RHpGEUsTmKUWztDmnmPjttCWSv5StkEqEAfGK
EUFMGPkXIaDPPlu4tKcr01zih8KpZ2zT71e7lqgQw8dovqXQMAFUBruqid9Tmz8/MIwQyvlF1m7s
YprtjpmsWquAFQ18fNmtTQ6nwwbg9CXWBGQHSCneWdEtrEMZ6jLyumDT87D5hoTbwHO8XYCKLJ6Y
Pcx8QYcdbM53spHwRqjgVSv8OR1ojZKSAsdyKSk8pnOJnS8omD9LoxVho4IQDv0ILlzNiJJeiJh3
wzUZaLt+JaoAxKmDXx+jZp2lxTujxwFfxzKuD/YtJCbOnZKTizMW43SKLz/uA4+LkyO0rm75vAkV
qNlagYqgTDugsfCxHoTkkEUoVqpPFj7s2fdMYrSBiLIYsU7z6mxACCWAsbWzNY64P5fjGpGGzu1k
nv1GDEGkigzEzuhOSAqK1DwYeruiYsX7SLkNYtv8UyATy07w396/O3XwDfbeNj2zuTQ3E9vEfNsg
nSq4IR7txM/S1OvEecPJ7WgrE0zoGRJhSdLckm9zhGvYXiRAmoN9tO7sL9s0YOPMdXZOstqw7xQV
QiQJPmhdrMiVqXSzQKwqdIAY+tXaUQyOkd7gBmCTtmMDB8qEPLla/jS/bdQdOIbHFr8wwAQMWxwP
X8XN1Pm/CPWgqL5pRpE2WytNIY5e/B/wLADvnk55gVRn0pVEkTCzFzo9xj3mKZMcBLZMQ3nzsGpP
GnfoBYfFoEKN9ihJ0glYmPpLj9KQf5iSUc+AY5SbmHDh/uDPzdM+6fNYYWarfENvjHbFM8gydIk7
TgOUpHp5AGRkUff9DwTTo7Gq5KKmZ4M3E8MiYdFZF0jTgIo78rkkxh/NbSQbw2v57LSGwXvDWaC7
EDC9AVTv+wHyswx5paEK9B5jka2UT5FtJy9QPJsQrUYDtJtzSVd8XqYLVCEavx03yL4651KPcA6U
CBRC4xF9rIeDd+DQHzYsH3WOcYXfFvagdie5xnGIb1AyCgGNBUU7ZqzS40IgZFnfUyH0wUjmDSKs
AQ7fKOe1i776HgO9MxFoCoAdrlzPeoSuhPB2iEsA/BUxixHb5k7UedL2ba1diwC00Z8vWSwMGX6g
91IZIg7oWhcWqg0QUvToBeVOIFh5SjEw4ek2Vd3wJPH3d2Z8/sPu9wkOJtT1iZh4vGoWWbJzLhKk
X7yU3NiraUBrKryKzCW4bPbcmWUqfJ7igzKOFhYeDKGyYVle9vD207IXm/P6yWuo1nlw8tYEnqu3
pLBEIwL3ceWxspcmqlP4IIooxi7ekQNdVppj4dqefoEENIDXYyX8lD5JvXt2DllRSGEUU1kfkUPX
KYdi82F8aDHesJ6XYF+6g+kW2HzKrQmCcrG5LDZvKwLvBj7p2DHbjqxf4eIn/9wd3+lrjB5aUeY4
dcbjRhkGEEbST7drUQuqhNQxopsQO6gHQNxrOvzwGOorInLQCVQxkV0sFlUYxj44zps2thdr0cHy
LlEnqXgrsXVB/0o9VcnGqnwWVD73301u6MPs+jtu6O/+0Ge6lcVzPsQSxfLTnTSJnCn5k5a+nGxu
C+9Cg7CEa7HaSGzWJUVbZ41Jf+UXMJSqFr9JGmLJTvHGbMQ/qMR1ZTEElCB4avACzNhI6fyQmI/+
1Ue8hrWB3Smfkx6vwY8oHf1TzarYZtxQK4dqdF2yZ6AIchIQi9l2b41MKo/MyJzqDDHwtpL36pYF
7Yh7kU0pvycdE2Gl6xWRp+9D70IgV8i/lAGuMCmq5suyk83dHRciQDwnDPjgCHJCbjerGgvPuYdB
ZF8TbOktClRpl8cj9auZlEAmOKs3EKpHKPpeaBatFRSS5ZD/elUMq7lH3T16glPxfhC79NqXPTUE
a5m2aydr8qBy7eIixrbjV2XEkiqz87WAS9/PomdZfem4h/XVwpmbGZ3TWCqsytfxYVFrjxX+Mnhl
lj403ipk/e8QaGbrqjOw14dr8eZKfnYS+JWHJeVoXBOw29WFdTl0ZlgI55iDaITw26q65Ztdy6bB
BaXLv4HhwmZhxNee20kP9qsySa84qBSP0FgeFRFiRix3daa8z0mvyzxXkwezNEs2NLfj+7Uzg54A
4XVk6mHgiwz3RnQRtHB3dwKyYzjfpgLUalKFHdiSB5H1/F/BSqYJ7dB8nR9dfAoL0pvy+HrSKdYA
8lB7R7h8sBVnHcuHl9TZCH6Wng/krwt6U7nrb1hM0QKqb6jAs674mHVfe6+KQU0OxXhhhy1mO1+5
DnwIcVq4+QA/DjP4ExivEoJaPA/JDcKgbQB+9sCToAsxima8CRB9EeuP8BqKOS+o4pl6WxgMWr4y
+EGo8WSwUvaysIYXEOROJ9DxsJziRQLxTXSyhGd22PBQtCGJFNpUo2KyynCmuQ4GJ4LNIVG5TkPM
P7zi0i6Fu3CfO8sD5gYtpdWGHHmbEqCkomm4j7BfNPgQdCAmv7hcchX5/Z4DWmArCEscTvHaKSCE
4yPA5mHtI4nIuWlqYwaen5s/PUDQZZD6b3PNdHU1Cf+NJYpldFzKWzW5DzIu/9H08AqdGewmqh9X
dWwC0b7qUSPRajdZjKQ6maXXs9Fk8vA6lnzkTPFZo6pfrUGGTloE83iUxQUFp/AsK9tTWaFIkQND
w0ixmy6qKsP4JSMFDfXdJaO1n1ZXjeF1i7ebYc3T/5w4MVG7zMyNdNU6XbyitVj6e3wOSBQn6Yja
YOZsK0X4p/Ej5sLJkbpWClSRxWAKR5lUl9mJpByTmiieaRqqqcP7iUBelAYcFe//UAq/hy/29wy9
UkiiTectn6CzP/iDjBxwebSXRYPArQ7qEe+WtpXczQueKEKHPmtMoHXXnEa8UjGZzrisRTPtdIjt
RyimSwAxWI4BmFWOXn+EcUs0zXonE4B16dhESvBei5tfWjL1h7B6mUkbcj/b6lxyq+Urr8Y6NJC3
XtsWYKi9o1PFLyHzK0+fgjmLWJTte7soq6ewZ6hswYA71izWxKiEK+/Thtt04G9wJH6cfBeyv2Hk
sS06CQDe94n209wMG1DdcYdTDdm2mgdQLIJ2C/nM5GFsgwHqtBgrEMkCfBI8bdws8Tgft08TKqf9
Q3Cv1PbXLoREZneSELY0BZCMjkhneClRLYsRwRamOBKwloMcHi30VduKl6uug8W2XaYxtd4VJN4C
KHpxwpBThwckFiG2isqNy1gOeP+F/CGlHsl2jX6dAOJKD4VUmZDsiYGejGMNPn+8KcPRWHkZWLk1
KSsi93cT5AQGA1nyF+SSzHtrBxwAKy/h33ADWwNaA/KtJLGAi2h7379vzNFgby2RDN9qB7soaojZ
a4T0aNDKsr53XJjevf9ZwwfE1cta5v3ZFhyuehX+g0wjI0kjfz/YsUzyJy6m/bn6msHKKmDMN/E2
EsYxRhDJHcbmbZQXeqecVelOpkqzu4ze4ZnfyR6QXeAu9lT+miSK0kQmW/RirA82+w28lz5IU3VV
fZ48QJcwqwpklFJougFNHDzNcnkBfB6S27xis9F+xjtDhJmbte+3kiK9CU6kKDC1VQ9EeqoocOWy
Dck2Do3zscuTIxH3AD2nCLid9+mfMr/Ib+WRBCZ9HGy09UUgljm+EDukBEHrmRUEPtDHmV0X+tj1
og0RA/ZVJstT4PBfR1D5PdRPkMbl9IRmxF2S0t4S/oXoy7V6B4IMuBEb0SWcQP2n65U+jDuQxBpU
lULEL97eXrIEfwrTrNvDxEYjjMt3+UT4h2bvPrVp6CZjp5DBDfaxouX/RfPaYNfmv8V/yLLqH/lV
bQxYssMXmA2QxqH3Nb57KujS9J9HaFLzRr6pb/yIdfgm+z2Ea4jyU2vj7xtYUsM2p06ObMJDr/0I
PuY4raHyy9pRiEfMWPxTppjA/Pi4mwKrMKTGk13PnpPrBojtnLNFmARriT1GGlwnlaD7uEsGJ7a1
S/VRMKKoa0uLq48r5F/1HQw9blCMAizhy/cq81jyIc2DDMinOEnhKXb14PV1Wl6MWS8CZ12jVVKS
JUVTFIAz5VM1X7xMo3ywfhg6h2CkMql+durMRpj+JnK95eSfXHtpu8yheVhy/+56ZeY9C2zKPDMW
xP+ih/J5qtxEipjlkUSGgANv8MIw0ijIeeuvNNaMtaU+S84kS6yReF2PSLrz5Ec5FgNz4bvAhGTB
ucecOp+qUso1ClAsSU9+KUN57m74QVEe8D8jZ3ftQX93phZpMetM3Z1NaOjySIWIXlSq3kh3PM+V
WPHwouCss6AGSG2QnMuijDbDmMZ0BG2FH/4KrnqrjiNZyV1pYwljfK3dhQQBcoltF0tdy/vSmuEb
vonR5o61GSkUwcEqdCLeZIJNsNUI57YZguehNuzCgkuR8NenEMiXQNbSXXP2qVZyKiOeO6unKKE9
L44v92S7LCfbIn6KtPfPa8+erTaAy3mnHOMpbZk+UninVVDcX4AUCkO1SL1czfmd+MLntkP4nmip
vUyC2OSJf9P8NgA9Geac/9kERH5YufiD/JG+dyUoLzaZtohVB13jdEeU5zJm9pPuen3hVXpgVPKa
BBxS5+6Xi7lG3F6E8yENaenzctFW9Ii+1FaojrvvkTofPbOeYqN/BQv+hkAumlPeTfEol945yBCp
o6HIWr3ouD/DEaD6fNlfV21maUboPQhTXikMSDxV/kboE13LSuzDA4b9+Sh1qeij1NsYCqafVw8h
kQeexziBXVVxs56UN9szr/cTa7WNM2jfiwO7Y3U6Agpcrg8CrSzVtNlARAXmyfQCgD5QD4+dXGf4
1F0RTzfcVD5BntqC3K2WxjFqk08DIyIbAg0r8BO1kVERpR2RBh13/Af4HSW/nVLHSG71xrD+Dwhq
Ro8q1lZWN4YXZXwaVH0yvlgriBU7aDORs1zludG84jlaTSL2/fsYUC1vLtxBJByxnkyIHi21Ay60
LcQwAIfVFp6Drz6WRpPytKzb4wgZOyqQaTdHpCBHtD2E06MZsusJtYAxXwkIHENi66HOqQ7YM3dW
OytMgN1k5w7JVOhf7mglM677mmX6sREgsoLT7HMppVCNcB9cI4THN8E6c/+xMJhRXh5yoSGES5U2
SsdT8DYsJRH6L//gZKtFpwAE9MxPJfwamOAb16zjJrVVMUQ8KiucqCDoocqmYqMD8JgZZbb9RinX
F00Kf1UsDqRfnkaxqBECACdE4z7AzJgCBZCy6lPMzh0D9CYh60/NZo6S2nf+NGr5aPcZ/u0PRzKK
NZmMjJYfTbGUID2EKG+MGgRcpdn+jo6VMvdDkqZmHSazFK5x2QqtN4x5PsdKpind8tSOlzIJcVcS
/6h4ASIgtF9HJ/qGXmNjWpyEYEC9QMTBx6D51WdEJP5Jk2nzwUYhWhvsijPbW+HeA8u5o6uWZ9KF
jhHSqsSP2LQz9SBZVzMwgd6027yvCP5y2h1Ukae+J164Pcy3NSLO6WaNGawM3Q/A6xPCteYGGATv
nJ02V2EIs9RBa71YAbhLvuyZ7ziG38bLhHQduO0O9JxQW9zBR8bcARufYRw9ikfGW7YM4sepAVh+
+s7tlAkMsUjEq8HtgACf1jA24wKqpW8RjUwu/9cB8f971//kmtuGP/I3pZjyh1Hol7ZljQdx6SY1
rfw2vpXJNxIS/9C2r0Ofotjmypy8bpePnOocnQhT5ps7pspVrIcxh8NJJkidwbIWmJFT4vEIvM0K
SDzPUy3E1PDl3wsvJuwQF0WdP87nFaVcnBwn+NOJE7RdGDfDFusL6IGczlJtv4F+3TNCLVyLDIXx
+FIfiA8MaPVySC6piCKUE2yASmgzjVvpciQ58PRMk/mE0244gC1yGmRqDs7uSYvYT5hO+OwieEm+
15kRsEID1fZzjypfcKUUUQD+frltESffhznS7FK81sLb/hKsd0PsJL7GJ9dJcL/Z4T5T7OU6S4K7
Svy1X8zOvmQA0LFyYPfLCMvfQSLWjXBYLY+STgLMK1uSD14LBvcuYvymYEdulAJpF/NyUJyGwW6M
4jWmy5F2b/E+M7ttNNmuPz8AP58edXxdMG8cliIMwcfNx24cIbtW7GQjr/+REQJ5VIuh0VO//fVB
KKLlMeNOGxbWVkGFFwul7uj9zeqbequ0AybcCsQavVhoRX62CvnuLmckP9C+MCmgInGpT6PEqOnV
a+XyCH5sZyqggKgTgmsK76eQmd3talH30CL1NBvlu6c/otsQg8lKKjNGdvyynptvuoZWDxAH8EKy
jGsYEhrAn5PxuXkOWo7rkQorJJHGg5N85p6w+XKc3fKOLfYwwmywDpP5rc3drhVLb9PmBA+R42YO
j94+F/lJIjKh8VU1TEFWfAwYsaFuwUuy6tV+hqTMinLR9GCeWZHnEUzpa9xi+y5BiXQShZJtHHCS
wTh+oX+xK2fYqp82kwFFCqO4bL+CmnfA69Y97trML66Y+D9c2VZtO4muGXtZnvyC29+lNysT769G
QzxS0KSk8BCCWC4CnJQOGherXDWzQeqjUZlYwm1iUFEz5cNgBPfccRbSgs1LzjbxO1OMn25WLp0j
JPqQ89B3P5JwM593nyoXm6T8yjpBDH5zkNVXTAmytKEuKWvs6/JhS4J/TK7tuVcj7L7bnylwP3H7
Oi0UYht4HghAuCkq2AFKeKHNEDzs9+S/MbOZnaY+bvTCbnQcEuGtpHuF6kTDT0NOaBNBx8hMuVSZ
aut2MDXFw2H/yrW9zor4vKh/O0wMRlTYeYrTyTipYz0Bqq0soze9CMmXBbQUxWkaLtuapkxvQAVX
VcmwATitE8OSOTP5IDXY4DfLL8cqB8ToQvrO5zNpfdHu/3sP9yvMMA3IVv4Le0MKykNEaSIUmc0/
Yc6qPJZL4nCA6IozDDEVzjJ4qvhl2icuaKuh2tK54ZKa4qmCh6dR14xBtTBMVzlayK4xz0kcO3A4
/VgIeDiXwjQuawj3OWEl0EccvhJstHnMhZ7tI+otohdfhiN7d9EJ5kB+g4u0BZ3FnZc+GIm5GPG8
wQwET4ldDFSEZLTu7O9v/0+Tp4uCrQ2TO+OiLYT1ixCD3NnUPsnlEh0hc1m4qTqEag2TxL4b+t4p
jcmrL6/5smrE/cZJ8V5cb3+WQ0Exy+jKYu7b54BEi3aZ8xjATdJV6rLhWX994R+i+ntyHw3d3J6q
8xEiOrxyV4zscz8ecXrcTXPJ4JgthfvxP4/xe4AXy6HeLsHibAdPtrlyunZlKTN/jeFdtEKrBNpe
1DZigxRuJDMJ9+EuKucO7HVSISC0vWz8zbTXY+fH1qsEijbfHwM1545/7jPeTIJ1p9qYQoOo8gkn
SPO5TZ1wLtgQ/cP0Fip8bBZoiITy+/I5wDuoV9RtKjsezNWwf9YJdlxBaWK52hVMG4SmjVVf+Ov/
iDWVA253IOuJ6D05ROhnM+VOYwp/8FltXDPE+pNHW44r+7fj77r2AWSg+N2bIqWZ2fEvTtDE0A8N
38z8NMGmTbumM5vB7fvvJkJjBs02jnhmvgo5fXEXsyW7Rvbq2waFM8alMeec6MmwyevN6V0h5hrJ
9U1D6aBIhrpDvnR/4o/4eAXot722aDPop6JEnxbZcKyfRDCaBGhDVcaz/ypjBHaCSHnNfXmC4lYw
JY7d0/EPZRsCKDf1KX080VDT1X07tpPceP2TiS8C3aI8+oXH5kCEhG3Tc6dq3vf3IRc6IX8mlpx/
MsGxUZqG53tAj7cmV1cXFsy2CclWepEySv+4TdJrwbxC184C62sQWtfLYhlqpZpIuFVftTnJ2fuz
h9IbNOqS1+518gdeHEplffv7lbLxDDJybdoX4bBGyMCzHaI3vzLpa7jasGP9Rnin+fV2Rct9cW4T
1K2y6FvRff0jGUQw+FJpbQMV5KCMWQT1lgn7y0cAHik+86vhQEVXu6Y4aMzbpkfDzi3xJcT0JjsF
MHtKa41+yqk7ZszrGjhI7I6sKZyrGxi//MJos/pOHK8XV/9mgWY/I38sUbhjqrY37YWqJfqLE41E
HwwdwTKDehZxRUmlXorJDpIlwY7Tmf7ohAGHV1V3es4ixfQqfX03z5izBWCEu5S6sCyaUI2Sf/fJ
NkjnBiZkn+oOK/YxE7cOruGaOTMmvbEXjgLhFM+B/DkO9NMV8K2R7kuZ7RBkWLejbIy/Ca8XhcPT
daice15h8coh4OBHC0aFa5zxY3P6PehjZy06D4POV8vJxtRdNa1PIuUWByQgDqUindgjydnKkQrF
JGdo7MoDhodFbSobQKPJQseny3UoGDfcX8V4gd+/PMqdokGUvpYs14Nl2KY448yOVY/olB1KW4U9
3CfqCqGG+eyo/GHiVdwkOXhthQPtbVr0w31bVmKNr6IOVV7AexwpkdDtpD9qX7hJoz8d4wafVmJ+
sM9+xwxDk+Ee9mSG8rbyR37usxppuKOzwCpjEvrSz+gpa/5IktORE1/Cbbf80a20VRE3XmxyzbpN
eUXt67Ugp9MY49ewqFoPCBxOQ5rFq1TIUqMoRG8sQ70S0yc6H1qmyGPllIWBEwOxhi+voPxFNl33
YwH23AfJwd7OSeHAnQLWWGZ4pdxgJo4T5wR/SYCJmP+8cVsRl0bKaCPot9R/QoEtkANyLN9WHrST
w2co0R0NWMqKHIr64hRswjYG3R8SAFcEjSqJ82GhVm1+utGLAaM/+2whCy+jpb9MnR3DtpBk/eyW
lZFTFh1u5fkdXb0ocsrPZ6S79JEs2UlOJIhV3lDwHvkpxCPS5TwngorIrlZGnVVH/ch0NhhgWLL9
SVJS71cLfXt283wI1njtonAlGZsk3ZTFbUD5nIGMAZvjv0tTJqDYAQhmBo8BxLVVeH8ZfPgBZFtK
RqTNoWXORkuoKqh9C3CmHQ7JFspUxEae26JLchefKkI7b9ZIFGO1rAy/b5dREC/uX1qKf45OJazS
6rZ2DcmZlnVMCJCKcmGGYgwkELYewXOlSADfOQUIRf0KywcYLlYpJ5qXSbgIO11/SEXhH2TcysdR
pNtb34ngqo7cxHeumH1WZaqn5SwmcBwvIUuSm0VEk1HicFPU/MFKNgMicEaDh52rnX75H9IhUFb3
EMiO0LfWbEmHRVJULbg0yRvH/jNULjlqtD/zO7Xcpx0pNPW6BpK0pf+TWVeLQZ5mrUgZUI1Mqeft
qrGAmcPpdWC9CY1ea25dncnQbgbdOjC6DZzmSqoq5Q1jkJ8csw5boL/oir7vtocb43ge8uwDWNJ3
EWoMmPgNgNXe1BdI+0G94S+1FywD+/NaoejFgcW34AYoABBx2x0jChvFz3co0jGEgWas8sFxmz5y
YHoL+XiXjcbYgxO2BoCQBTEqcGHcKR48eR4+54w2Blhl8j/sUGvNb0MV12E9c2j7ih6lPPaO0eC5
NTEhDFvvcFLYuZZsuL3987ggsAKanPZekQEjUHCdnGTMgAUT6oHqFXTmugJV0/2c6AQ46i5zl2tK
AlX1hFAuI3O/ByYmHfj3sqiSS3gOEMnhGTG5i+US06bDGaa03GaIEbIS7dLFAv7HkQFFqIOmdmSw
z1Pgk2+4gfJfhNKerR721VeFUhLroIKYIglcIxrstwc0iQCG/w39/xTu6XRntW+Bdin3y24MnyS9
w8vTXicYL560OSNggl/PIN4yPGY8pha8iQno2ZfB6k3SmAYBXU2potaY3MlpI9/OO2Av2i6j73i7
BWqNtl/ERQ0KXzJnIX16Qib3L8PCo9GiiLxq+zDTDptUUhOzwNxLNLCWExioTuKmh9qEiOBs6paA
ANQN1VqdZwRiINlKC6BjyUpNFSH+tb6HB9UqAla642zlHIz841Q4pqYC/NM8ixY2IPRxkNdWWKjf
akgJpXu9lR5oHD30FnEMxsTwK48vbvpvpGHbjihqV67/SpMVY3nGhfgdBb5myD0PButFtWUknLe8
NQ6DXR0c584SA4xRIc8vw34hYh4jf/Dn5E6pC1kUDhcUZu6+FzahbEMEPwp9ck624TM2/xhjkbNY
r4OXq1WqizH+Ryo7dxZz6ZbnJcpYtwUW9EAR7oaP3z9TBG1xcYuZfHBjsZipP6H9XoCuCJMbo5hA
GpNyE+KYv2+QXDXPkvPloBUZ/z84Uc1CEviF5T/Z5DTKutqZW7BW/0nE979mqlo1Jvyknlp0I2sF
iFTTb71iFk0AqnfAnd4uzVpqdCEqbfvTz/dmVlEvo3wKp6vb3yNTa7KEpTy7b7QvrASv1eQf58Y4
OMGNFCypSP4aV4XkZ7uy6YWst/kFBm+ag0KLz3JZXA8PyTj/mSsvUReylcxa2jGZ+MbsG+mrM9if
lT29OLl4uXqDS5cVDgSLIMtin3Lm7x69F21vN/I3mbvnhT1WHTIvTrup6dU6XQtVmq00T5EqZS0w
4vt++x5/D8m862+NeUoZLVLrDQI5SkScL62GSlyzRT1OUgQBXRM4oLpmdYew82WTtDIcXfNHoKhG
pMyny7QZ6nfp4k0Dl3FUaMaokOT3ta05M3fKiEVvmcZy0YpJRMGxXplOS32XRNEQsbC/F42NVC+S
uQiEZ3Mj/TcEH8F6OwuxJIZTEhXirNjbE+h/wM8D/t/3DyoJI2307EQTWznjssg49iMJnukQBSqP
lsE39OEPys5f7pPlH6Qs1xysy9ZZzvDOq50zCypC3D2vknkQt81cY6fPt51UzhglJLLixIUJVJpu
PuvqPmcXCq8FsihITdikHHEG5fvCqOxKG0GD0OPtrjQnUSHokeiVpUQLt30cKjiHxgF9eGCJtCip
kKjuPM2PAxmaxYnzLwOYdpsoYP++CRVr71dMbWTaEcGEjik4bHUpppHIZX9QMKU6XT7l8g/rjzvW
TwJWTKSD+hGKrb7AMLtiPRT9ylmMhfF4zVW+2gXtX/myOzE61dArrcukxFZlgnpdEz3zE6gyM/2g
H5B/WiVNMV9LK3b7zs58mRL+1svF2HA5a71Oh4nwPQIvFZVa0l0CyxEi8Z0Erf7x0k8CGpMBygXY
MqrEiWjUim+I/Z+Hj2NqIApL4F94OFJwcbEtIQlqJ/roee2PY5jH4ixNkdBxZdQ7cyyMPSvgFfAO
McMA20QvDsJP8Ru6EgH1Y02AJnXjtQX9IYtpr7pseW85mH/D/BUyOeWUcCtY7QdVckez9/i/NHZ6
eVLQ3Rvj5I+obofdf2mST2OHHUEyj0DXa+JekbBj9GEp6WEeHK/4uyeCa5qZ3jMAuku4XbGEmRXE
yOtcJvvO/PoM4HqXzuxLDdLgs+4o25D/dzOJgODLSk18Cwr50oOiY8DBjDBMATSIpDfhnWo4hClJ
DWj//7WkBm8AOt7HdA/snGr0BgGI3WocoZUJEh4hm37F6uaSHUcQOzSqN1K7f9LZ5HhVamxTCP56
ju4zlmnU2cV863dJaLRB9Hb+NSr8GVA2DtXSeAxJyA2ym5MSh4Jo86qtIkI5iZyI+X/f5MgDib4B
EqK2pCFsOlKD79z9VKaFwfnnp0QBzb2hYhiaEoXMHDRAixAychQHqVMmKKrlylrEM9D6IybqMBps
8bTWOHBIl2G468bzg9tVs4kIaW2/SSzW2Yfok7SDDcHFL+WK4IwOTk46g0sL4c6Zsxn7rpBeI3Y1
PCXEGke1NeQM4RyFGRyzFn8AVGZY+S7js0+KSrRspAc4Iy3qLmjHmhDjr2cotb8ihfaewtTe8cRW
GyFAjm+lJbwAeUD6gUuujRFM4VNKr6hLa3QTGSCMDvP5P1T3ZmjESs+DUWoF29t4XwUY7gCw3Se0
18XW+xXUDNHUSx5PlolW3wWShjlBT+GX3J5bJthsDtsUC0zyYKWQUsjs/3LHxNlK8aDk70oe+Tdp
ExcMb/4EuHbC1gvpRBWa9SI/mHnTnQfvE/x58G8JE+8yRVrK4DBNgbg4M7JwNiwzntnfiKsD+OKO
qWyLohZXBKoniRDfqrL/u4seIDnuPXgkNoM5bVQigaloOonw3zTma8D6xST4FKvwMArJcoyi7RrO
UGTzEXUnnSFYsMjTTexBGhm9xJPQ7KrqyjJnAbA5x86oMc3mSpPMfPjpNA5d/EEEbawNhzvkX2O4
Vq9610Vm81M0irkKewvMuHFS7gG7TMWOQOgMXLjKxyzNIlt3FTjaFoN7WM07uiavNebiavUi6JVh
zteujd1Dlz10Ddt6PnizA085yVKOYwMCgYYU/MvTHCYBwpAxvhA4HNWl00Vv3DYO/KGOUIIqEIu3
LHWFtrZAlVtvsR2bkXlxQZUVsHbUkKlvdfuMZxWH79GTdw2R0No9uWxYI9firl3PorYZp7o/Hahs
MAV2W+RYAXBTT7dU0wBYOFBQQkVAWf2Iu+BvupKVxhpHOUOReldnLpSgu42Xy2CCkP/G78fJo+x1
JMsxkQk9ETAeq2acoz5GKXWU93AyicD/WLUzXkoO3CT3InE+ejY9a5oiVISSFoEnWH9NzttusyVU
gShi4covrTJ7dnxgEkmS0qkw/i8RSbZ1wZQTJYGxrPmqXcA0l9RydZbyL3iUJXpUEx0TYG/DVVcL
MDtIFaeU/i6wHJRBl5JNSuEKfQeN8GalgpHaDpTnHaUeu2haFvlR/tpAKGdCyy7n9FABGSQ0DGsb
x/4gr7qsWjjfcmgWum7Oanlxe8oub97zseeDqPki+xcVLp6Ms7verUNSUtuy/xVugkcRQK5LlpNj
yqBzMLwguaTP11RAlUJvtv88Vr8fuBIUH1q7z8IVehT8Wo5E/v8LReHCj4eaDWQKec93++7W54or
2gbXNLYDwGE9UPtD65q18Js1b5rIrP9uZClADoziz2y1kDTtPRTAroWHfbN+C0Kqnrj9TDTy7yvk
ADbfsH5xfqUnhWC7t8nFxLabHuYDp2qV/dVb60CLhv12XtzRfqHg3X3JTo43mfZqeUu/VePt7J2K
daZWWmfwD1VQDJ+3hfHNU/Ug1RF3mIdhZ+ajXlGzi43koTQCIwwwA0ldAS6PPit9wouNehWVl9xh
MA3BEjWjwzkS5/AT1DBC+ekLz9sIqbCFWX3Slc41QmV6G96YFRQv0MteFS8p1IqOEaQcdyX1dZ/G
/55wJIFnvqhtlXIOAb0Xum1qOExJQIwRo9tA81gvla/1Zfce1gr2wgBnnM8a4QDIcfzcONGOaik7
vxo8ERf6dL84M1nww2vHPgi5J/nKztRHsGDY7PwO6qu7ZZDN1Kb8PTTee4gkPyl21aC7wRAhh3tu
dQs4ZgLXCP8r7UCjlJdEt64TGjkMomYnuSi0kZVQ8Hul51wMi/6MR3aIwTYWCZ6Fl5CkY3COzYZ9
i4puLgO7pNvkk1ntEzwS1DikRqv/LATNLWHY8qhgfxaUrl8Beml5VDZAnG/hdknxrhYDzOQzaM4r
Uphl5QlPkXt/tsS+MckINgJSjIYLeLESNNb7aUEeyZmuGZKRDuEObg6ErJpbdUuZeh25N+DhH+9j
bU4Af8KF16nGDHsJBwA1q7HLziufVu2ZIuFzBtN9+Fhx9+b5fApZskfn3n/URIw65JxESBagnz8b
t6rTvWJePhxKeTpjRITrImmGS0xLSEEtn28BHswkgf/e9WjyM+uhic77W3/Wzp3f9/Avyln5XsLs
mXLJPT2Zf3qlR/GW+d+gAXkEWTx07w7Fo4fpye8zImbjkIy6p1+zKoO8pV//IaWviy0Oz4K0ToGS
Dms62RB3+Alm8lpLUNP3X5Vd2ma0WxMeyyV5BMBxkK+96kUMkhs/uPldfcy+huSmbebwUQ6HEC/b
QPPoJCGTq5bhhKyNOcKjj/3fMyLHm8Mw5SeTSXiAjeMZ3DDLdzNpIjo9SNP4oXpY+4HaI4nyFnzV
O1KyR/6CNpM3rnPDqO79dOEuGz73KuVQvz75ti35wlDnQcU5Cc0thc1x7lIdJpKhM7A7ghCsGvWk
sQgKPJjcQNU/djYhDZBy7km5w+N08akB7ANfYoo+kwgTR/Io8tu6d4b+Sxkz/n7nYvgR6nwRSjH6
8p/xUtEy7rIEA5Nczg9vpNeeoTrzSnCQFiusOKHRGFldwHj/c1SksEb28dACn3+gGHSdfNIQQpaz
jHUUhbsQtLnY2uEsIbOVNCdox2P67g4HhN5loSDIJv/jEmCfOJUjVJXm/qG731uIVBV6EvLJZ7J2
hcPoEEHMJh0JbxLal2ZAanLR0GsgXJ6TCUK+L9br882dbadZ3JbLZRSWI6I2GHHV2d81AbewyaPE
PMkMZB4G96T0ktCjIdNxQVSjLJ9KGsLKWERJk4G7plTnRl0RyF4uvyCj7OpIOYB0I8cqErGNez0c
h6bh1C0ILettp0jmIl+1IyIqpvddXPooAaNCkoauJLnUekfzRxp6N7UXlLKHd72NpGaD8PhR+tJA
D7KK5L9DybbEBv1BeWeJaud1CWMHEXASOlJnPVwmaDux05DVwL3nENyQHrew0SmCVzCXsYRI4cif
avxR4wn803OFa7/TMXdQ39WLNnvH0NqSH7cuN8w46jWNlm2lrF3gI8DP92Qo0dIiYSiYAfF6vpUY
jYfx3CgEqcLAXbIwzFcTYXHpIBWuOsIFyb2b1MlVR9D708kxUiG2cheVh47EiOLMXEbxxlG5mfG1
YVcalzcS89p8jDvH6tQQItVWZnFIom/6/OyTNP/iLVFAHrZ/ySAKv1pXP4U+FC3nBUf0UeikSQ4y
oR0NZz0Qsn6J87i2mp41y261jmj9Uo59GNi143YMUhAQP8MV7rfZabscShBJBEm1NhCVCFvZSMsv
R+m/u7ROZ2bb593bVKe/MznTwabdC0TURkQh8+4/41KmgBv+p7CWuV38GloqZvM2G780jWdDYCLF
CJ5Coxhd/fi21HVNa+ELK1bd1UQEKMcNWVZyXJMmj/oXb7C55t4j0KNpqQKsck4r7vwEmaw0yL59
peW25pALorloaPeLT6RQMn2adudF8KIBslLhHy1BI/L/Dmaa1sBtuAC/3/tEOAa7bQ9/kIrnYZZx
EkL3jmAs2LwNXCjXXxGLBMLAd8jPACviGC5puHtaQjHT2MB8DRmPi0VJmJ+bE3ax9z5tZss7alPC
X7Ithi0xV3cGcXkovl/XP3zz+Q79h6nP7da/ru4pAYh6wKIbG2nEyEHaa77qwwKkHdAbMd2MaNGt
KreM5i3kI5+zr5cf8CuAglhkuS2TwbQ/ljhET4yCGTFFeQ5fTD8UjmKxT8lIxvQFUkSyejG6PSdv
Zoj8lZw0q7Zb5cMgvKZ4UEnsLwyG7B3mgBSV5y0OPEZsoDQblwA+fAukg99eM1pLBfGbhK9zVOuo
u0lRA2eNGomgKi+dLVCWI1M1xUuSFQyvb22ZBh+CavCKyvSVDuEQ3YcSZGJsFoHtnnkapfzD2XCW
ZjAHC9pzxD5qunCijDqgTvO2D0artmmWCjBZl3y+gWMS7HIFPj2O+uG0xQjhT0/dZ0RBhxSu4EMP
khbll2J4dRVJ3d0uMbM6ZOpMptjou2ABujiTCWsJhTbH2gtPGKnE3pkwbGezA6clz7mSbnoChYfo
KdnN50FtW6FlnnVk3gv+w2yLPcoiYWFtytkvdA32BDBNfwquaSTCqHrKwCvU+g0t7agHtTsd70+q
oRPsrXOfpSuDqFb0001YPhIg8mDdmogYue0iI12k1uojECfvtv80aiUNX9xuHhsGhCRDto3ZvzLS
85JEhsxpXdAMX56UAVdDMj7bjuCW/7ttID776v9ohlnMRQi4kf9gcm4UH8u5agcxa94ab7cIdimy
9ZIDnwJtqw7QLYcVmjC5NnClFlY4kZqZrBkKIQCK5o7o+B2Cz28e8jl+szqqRgyPc1yKcSPXcIS6
AqiTZFMWc4jNukXyymzmm6OiczWo9I/FEKVu2LwWEezhn34xQ4vBq6qjTu4wnuPDL+4LcBO9Fot1
ywNtQzHfiMkJ2efZnlQUowRxrnK/ViSLf8/xlRTbvpX6P2heQr8ywgMJlRcV+NlsqOx8u97xu/NM
079wSKlwaMisMZe9hAZHMNzVi9H4B55nFejYf/MWLSDOXdQBeML4SP0x7ynupP8sY1jhvQOQW12/
V6+QtUBLzI9gUxfl8VnkjrEpsvH4QW9IKWvV75oi36IuLCdllz7XP8cUzJApc5qfqpXzRvStxgpn
qSuLivkJ0EAZT4gcwKsS0M+c2dN7dVcmO+CqXsva6nNv4g1/t94UxWk9qe8536yf16mT2DXpTFgf
euHZSMzaII4M+HxaBMqDFEQwmg86IOxU3ObZetArK/MPsXbRHwPEU3AwyplSkgSbD1HS2Ne6XWpl
lDmDSZAlKJQWLE/ZAftazaImlUx9cviJGUHF5TjBi0p0vJdd+kYAkZSyxdqhiQFjxVko9LCAEIgY
A6aQJAeiy0AxSHQKGLtkzxkX+0jSxHBw8Yz7DcibtqO3Qh03xRl0RiS6LahfHSzzQn2k6r+RhidQ
TVVjDLbLwDTGM4xb3uH88piccGVetiOvyfy8EG3o9aACtrkFQYOY/tgDIA0xc1pZQtU1/BoKA7wl
RW4nEH9QCOm0bRY5Hu9c9byGTwxAGvJFV4VEGUIZdbhDzjdmUwmAl040l9GdEiJltHH3AnFtiKXq
5z2UFKNUKqEpEXsTvK7ulZ8PkbVi7jNIyUFp24yjwppZlgIVIVrBhviXoj2VJtNthmdB0vHEAhVc
jaXUCURxFFZczWX5S9e3TrbLPvEMeNgmoZRHffNP3uB2VbsZgPV/y/xgCP8xkYIXJebdHzBdeSDw
tWiJ5ekWOpTay5245Zt5VCEwHX6q6UEpXzKsRZaQUsIlO0B4dY9bJHtwdxUw8ydUbq60qgH7F29f
ivt/oI5yzCPQxWnsea3yluHdVF6UT17qTrE4fmihXGcT3oTXEnbm6xoOsIpqEsLcYQgYWl+h8uxE
ayYzfKQF6FgjlxlJCTE3Kt3BXZHdwnWI5kh+9iC+WsHZMg09O9qvNwUBzh7v4AGDQBolbz6Uvxpy
331Wra7X4LPM5WN2RFdIr58AhcvBj1vkdOn3kPsmG9Y4LosMkMV8e4q4UuGZFLBDWBO9pIHmEJ+W
YUrnPer5LPCfX37BdhyHPHPcH43lNDEVZcmcaERZvKgU8/s5vuI3CjhcCkxIQlSdcdDMbKE0XSeI
pRaGpMEykHGb8d0cB7Ji7DO4bgegUi75rlCtfo+FZub0TRHuEwewhJgT1q9VNb2Kz1BirXmfmRSO
yRvB7/Aqr+Y6Sn+SvklrTqnuZhaMEJpvoI/Z67OXIBwsmmUuVIojfc76Xj+CjLSDF/YnAulQ5kXb
Ewe2MYK3yuukJdrp2TEAKVL+LT0NfQObN0b8A3klBQgPDt76Owvu00sdeA5PuogDniTLHFYAu+5/
Zo8vJhCWYT4Q4LTT5Rv6MLF4aYFwkkX4yYkCezUoOUo4yRzu1wc0HrZnTaQRSnI75vst7W9SX3Xb
OsDapzo+5rAAxnGpPwzpvnb51F/lIFk0Wr6bB/g79AJdY2JDqiPk9nLH5TPeEzUkzJ5L7F/XMkpU
ylKPRUr9Q6vYkSXGHTQmjQVtqQj7AQNR7rPO4Vs77JuokConkJ0pblK7ZMFHdH452gHPyrUZwneg
rYexBmybR86Nks2S6Belup7wnd2yLGcx/qZ+wCwfouREyuF63Be3/pYEdiv5e6pe2vMXQ66GZiPp
V7PdcrI4lJprHkq5neqfm9zaXUg5YjpXSkbGk616GqCzDtFayF9rVRbl62JbhpfjsDFiVWQawiL/
QW6uUeK+mBdMhGwxPrzG8jSxEi0P439GdmVU7lLyCVIBKLv4d16yFoyEoqfvPUxyzULDkVItN7O9
PKb3VaSLbvtjH2O44cUdfg0/IYkCiffCz+x0H6wOWgS79hNddRhDcWKHcI57mM4RxQLjZem1xTZl
JcCfL/z23mRLHrNdk6yAqJUFaY8rL808JWa1atOJK6j2eqXJduNpnVrKcnNu5ySP1GvFL4FTg02g
VnG6yFvpQxRlp+JzLZqNN2rOYR9UW5mbaTT7O7XK9dAXur0MV7835VN/zsCM6fs0hAoYw2G84a9E
SGFDXJKbYCzeHaW9konCBIKOIa2vvrgw8NlatMmBDOrtk67Q2O0SNll5ZREmnqluEhKkTpFqb9hx
phaxjDGXRWZDuFg276e7BUHaVgHVcEnYVormyCCvjwfqdunHvQig2bu3moM2/wUKBRtCVBhrNA8m
02y+d9JkyIQh5FBt+GeLslAN6qlPoON8Jkbs0OhJcs2Ny9x2QY+r2/VM6uheamUQM2/aJmQevzPg
J/S5nbkhqxhzBZhKtirGP0/oXkwnyiBSijVz5HjhvgK0qDXK508kuigvOFOnj4D26n7y6tAMs1u1
B9kNcm2kIYmUAbyOpgu/TojpVoJ5TK8H2bNCSa3qWa24T5E3EHr7J8lTYbbUDAf4R12rTBHkdEP1
f3kQaduOHhb57wEF3iTdemHBhipxH21+EsxZmiGw0AlUr55qiqIEEiC85pvMGqTxBApkccCvzzWu
RXfvbjnUM/pDvodv7fZMp7Vh/9OF5LLqkPupD6mosUmFFMfMv1kR8dcUYzCj2/vrCxQ8AboGN4jh
IdKDsauWbjIErmL3TYNoM3J5ah/1TzdY7+8n/Mz6/tDIh4POxTg6S0TmSD+NGXg4uBviH6Al59JX
l9APvNGzmLz1ayDLJjoF3yiSNpQwiFWq5MSCfwSojedH+o27E/OEM0BIv56VX+2TCmM4sae/diQN
h/znWDV+xcYHpWqEHbjekoEOqMcW1C9Ul3QxmXF0w9qaUv5V3gVvgHmzZ09cLup68tOLfb/Lc101
hDvRF4ybwNifzkTHK9SzwjOkYM7Y8MosIgevVC9Tpm4NIH9oma5rYbNICmxw4Rbc9IHL0XO6yibD
Rr6kfFH+VSaEBiOIfNRa9yITL1psgnmPtrcgiWL00RsF/kYfZiBzHN8TXpVJTBCtHoHhFu4HxS5r
hh45SQLQFiZKBMfYrWuAhUSLvmx3uZQwFVoMAieNvUiBksLr7PyrlVxUo8HQIGxq8onBoi7dARVe
+m6DnWiCF0MtTCOEpOzSWB+pqFJI51ndE89IlU6L+B86ttLCv9FZSzwTB2K3yghtpq9acrdTiEnI
ybUABWE5LSwX7M+LrIQyg6b4I5kR20z+zoJHEiBs4GduH4iOM2iCZtFz+svnH8l3H5dJz7AIUEs0
5ybsxEFtgxuYs3tpNL/5gCOWpdqxroT4LQbCym1Ug0zRET619NwNuWWeNvSqPi546Bk629bx+3Zf
KEl3v/0ReehN0lJ2MVOp8dNMMhxCfJY63oh14MihEEhGLqgEGmz6zeDZcLB9apCQ9FJpipKhtlCN
z3ysUXC/kuX7qaKleG8Xx71eBXMswVSfsOuuWpOSNzX0iL1dmOBF+5r36uTxwZL8bropgQgxSwNn
GYZOhE0j/hi5GQUo0AGmqhfAoS5btr0UhRcNTLCmfz1dJNkdGjpsnjwm7NblOEfwvs1l4ivK9J1v
C2CeX7fS2pM8By6swoEU8tGYaF9KB7m7F+nYz+Roe6ZHN1/q28t3k4CLZAjo61/w+Ne5sTjzGGVg
a+nCv115QpsEdN/90g0VK/XBmEJpawILPzEDS3fSlont8UkYQRogACWW5ed2Hew8WTnrnkzxJLl1
15SC8JZHtl3wNIfc8LhgD98NyhFydq8vEjV6tjwPRefMzbt98SXhDcP9dyH8AuooIKMAxSXkMPNa
wiN05+Sp4JtFv752qGyxmvAkfzUuCfYaI/GPKIGaLcDxyyULXO0oNs4SCqkj/zf1f04zm9kGLqkt
CtIlq2W3aqkbstwd7nonq4pahPIQ5/UqBAxl0tdcp3Ta2QNE7RbK/MTxZ3iMWtvsof3Ko5+EZKa/
21u7q7W9T6yIMHAbx69YSF6WRJIWTWEo7kZwzhE7zCRtBlHL99DUqiGACUnXDmZ3fN8ZiI3GXHv3
9kfGoPlvThCDDupMACSJvMh2ujxNo1jOpne+11fJOavs/A5ok6S/0ZsjcZFXOwP6Qel2r2jBSURb
SiTShuJSwvkD3gkOhPn/D9D0SXv2/Knrq4X9rciuaUlgiCCrv5spaqQpKSFF3V9f4dV/wFMPHi31
+M18uKDOQmxJ40el4zVVm+lTcMv8PZOSRqXGLxeAd+0AHcANlQwSsTjOJkKXUugwaAqPesqubbBp
jE6Mpr0BwR5CGm9B3d6yDq+RSSfj1rsnd9hd3zWuU607ev/Xv+j5sQLBPYRIkLfRO27uV8QTH0u+
LQ5ebeWgR4qrfYdBvN1+VOq6U8cXGGDxbFWUtDjXT35g1H75MuxT2CZrLlvHY7uZ1uQ+gfBbUNGb
S7x58sci3Pkz5iwpyUPOGtEKJzWQXtRRNukLqn60H09sipe3gaodD4DOVgDfBK5n3ICoba4jSiwr
DoyB/4NRO0sEO9ZKHtwdR10ia48PtiQYl+W6pFZmHPYnc96DDqaZYelFlMGJz48U1jmjgYJvg+L5
b3CN2yYefnMfoES8yUT1/+29yOVooaEHh3uUWqfZh3Hmg3jwdjWQ+yh4+xQsoWy4Rdhgzr4ya1zG
GxrK+gX7r1m3W7/s4RTH91cquKfwSfpjoGE9jXXxmQjwqK3hLvVDBIRazoOFdd4okQ824PraRb50
gGo5mZNCuYPx9PIprNoVqzaqJ8uUpdEyXX64ArUChSNkjS7lknt2Pu1NG3STklnVkV4CGAbiwP+N
gT9nkVc1ky5dHs/eJR5flDZ7cr5JyN2tgdGBt/YGpvijTbcQwrQNkgqQt5C7Y7Kty2dRf6x9nddG
UZEamKNslFLWUpDXAMBq2cR08emCj9Zh4G+Y0CcQ2LkQXfqECFoOe1tKq251lE3ekVWNoOvViEjF
8kwSwHq0YrhDuIfT8xM0w+pXX2DxGuXJFRDcp0gTdQ5RqGQVFwUwE6pRuwetk4RmzuzfJIs+rFMN
qM0DZYKSHEoyz0zW3IJiRXlywFICR2g0Tmn77qaiS7WHIZ3BxnPctkXgpXptfiuZBDxiX9lWlxOV
6WjplOZffmJa04XkjbH89VA3dfb2lZcWez5R6Wu0a2PHgafKeAfUamtpI4ElxDV3LV0LDGcXAsCc
pkiK5QVrA45x2pFcfytxl4nUaP8wPALqyWDgM4VWalxzZi7BgQqBlGAHfIZL0Sxji0aVHlRIJyO0
yK9+ZsOilbCqrCRlpPY/sVFbPTMxaxcfiruOjfVXHoVvTtDQSCkIA5pJtiZS5Aw6KWG28ScM1T8e
Pb+aumK7m0Prz6flpORj5Yds0BuvAxrnPVb4BJmmimHF3caCbzg2Rw0ju5GVfamWLyjel3tnV1Rz
6WjHmHqT9qE1qBU17vxzRF0/HHnXqVflkM7Duwvbd4mdO/yNczTFb8TwA9NX/UiYh9qRumdwyhof
jcTPIaxROaqAxPkJPdpmK7pumO4knwX2fiz/rRHEaDs4ouW12xD/EUqSKAP2bCwGghhRnRsymbO+
hjlILyKcC+AqqGPe/xwCvJGxBS3RL/ouTkNELPyVDCjELx2CMmsZaUzljmPnM8/NXi85a6xyU/X9
9E93PRmZoZe6em1O2YN+tv/YVNm9pSuDg8+hY4HN0Uq6FEF98NH3byS0YThUdCyP6MwtdB9sJiB6
OCT/keKNh6Y3u6fmUkUbN4Q3R3tQS4w69vx8AP/HpY6U277mIBb3/OGJu4KENsHgW/E3dT2jzV8S
53yaXaNs8d7PleSszzN0RSbSoE+ElVoZEwK4m1g26Nvixo+1i8xoq/w2tfqj31oRRek6w7SU075o
Qb72Ho3+sWhQi6TneDfk4BQaN4yUv/+ntWRgz4Li6mD9ULRZ4dH6z1i/8R3+rpGuVajguDXnzGWY
CfYC1p524qU6c8Rmvzzhk1S5JOR+pm/PpXCXwR+I8WSKMsyuCE+fOXgrPmXAoFlX7cyG3HFyhcKF
/zx9y/oz3Lf86QGXYhdIK6pVcF12u+1Tbpbm6wSFotxxgYiq/kxjRfYJDAdpARb60h+TcJYOG7t7
XwwSydDXb0ciqc6tHtl9SMOxxPjUXkM9VOR+UetEwZDmnhogsNs21AYnfnmH2lDM/wJeiky+CpSB
73lVnQAQKJvk9jP+1ElOigM+vn8NupI32V1hwRqU7jx4t0EkJOndwk+CeO2rR20KPDRsfrIwM2EI
SmdDBOKPMF42LIw43j8kMnNyhvr6zcGajTSF/gDv9JvlsnlgcCg5WIBbsqc+SQXEa5z3QziI8/pE
I1WGyCl7HkvAj+o5rN9t1JIzsi/Dtxpe7lbGRYok0t70yPQvlKDJjj6Uwige1H3xoL4KzJ9iHOV5
mdzTCG8ZGv/B7V+v/uli2ma3e9Dx90CZWKsOJdSSS2E7gf4+bHzRHw10ZHnJRpONZsdDcbHaorZy
UtOObE1yscXedUwp8nzXSsKj/ZLUAsRXGcQ0xeC+0ZIpyAESTOZLpAkF9+S85ZowaHDRLju3WweY
ISbsM78Xvb+Sbg4ZqGBzRJeq4yMCcfYjy3TvNLS4+VtIm+pGouL5/afaEexcDmDZ/XxGauRHNqMw
LfV2o34LmhPPQZ3PxMVd9Pv1ehH4h4lMKHio9FNtGeAEy67yGGrY8eXC+wZVdDyTLOR61LlRfqIA
9uwjhPfcdLsn2H0L215I1QubKFauLsx3vY5aAOKr+TP2fGBfJAOSLcsZZkJdeu9XEZXL6USadfJJ
zSkPHug1J8Dn5mMqrCtO7VEvthVJ5OgK6tRz83LkLY9s+5dIXP2JN0lij7+5vQXZLR5he1bH3MPo
fmwv3mju1auyGyHFU+hyrJM1PVFPOf1+5NG1f52ASODbHYwchnqRx2SCuPADa2kqXBXxVwlKLQFt
p51Mj8c3JXd7JkjOcKyhcd/ftyHed/oPVdJlyiRal18Zn2YJf8ZqGcHKz/voo3aampO/rgA+O+Xr
RaDDeZG0ryII8p4M7wPRpW8J/qUYHiSpLAWIeHq8CKY66nqtj+TApYhqfbZDg/LokX2rl3Pe8J+C
Zvu0dmMvcHRBbEuaMcuDLMJtqZlMzCpLXrLPxav70ALEgRAnT38IAbAsLsWce6pFDUWtYPE3S6Yu
8OU/ljHx9ai8QivogAWMb45PFoYXI7M5nt4xZcy/Bnvu5m+hoI17bS9uWI+2ggV5CPf74FhQ6zDo
tRjjiwDTfkeZayLqEiZjgWYqnoALbhO541TseW2TkuK9C6sEe2sSCq8LjFZhbiIYAHOKlCBTbToo
6bYc1a8js7LIZflSt2TTsX9CcxjuymLfvv+PUoFwc4H+bkecQmX05n3qQGa5VGrjj4Kiti8rWmE2
+OvJOZQ+QswHk/lu6mh/1pqbvcuWjrQkMDkWr6cGBAUPvVppouw688O8C+06wXe8684ZBwCm5t/h
2r0SEQbyy8nNvMsQwOweYq/l3vbKkMJnfzejR4Ot3wNjeP6IRabWaCW5j2H5c1lBz8fMwt48XkyZ
Hxk+LTVYzac7ia8b3atQ1ckQ+Co1sJ2uMoFdqZkILhEbsaIXrPz/ajL4LsRJKXaXeH6ueiLxYsqB
N5e7b5jdsqKCbbaYxKK1p4c4BfizCZ7IYiREtShGwXMzMACourgB5n1nS3ZPujQ80yIVQ1hq7H0/
5Q4S5JUSpHZcV628V//QOwxPWFEuO2NzRREnDQdg2iq91Aq5nlVSJ7Wm7YhoRoxFYyh3FlcfxC9F
28Cpq1l6LK4FFdH4zoqYm7NnjlIN9F0JDyWCsw+5NGlNEOxTjNlmuSIZ23+2w8jjyZaXX9BmCO1F
w5TfHLY+kdpFpGcYZfqt6VnZKMrPmUTJYU21ANYyknPzUKaBJraCW+G/EMtL/R+QX8cTcfTnJWTa
AscB++EM1GO6b5xthxiQDcwTZVO1XNmce5wdkCEgJIeGFoDTvs+Sa3G7ACXrc85H773adbx3QG37
AZF/DnOUwro/jDF4xQRoTgXw1KdZLVdAd8BY/ZZeex3MORi3Sp2MFN8JDFzsAFKKPDEtgufeXowd
4QUECgiKCXbPMWLp/cq3KCrk4K0wRx7fjOEQgp3yx3BloSQv8wTu15mO245ckIlGIcKCTzTJxNIq
iwTJoGh5miWfCXwRFqPCv+lSH4XJ+jMM3O/FUeAZSHBS9hZnlJpycdeKAF9gtE3HwmT1zw4f8Y8/
b48zfRpUlntfhrRgNcr8OUTqUzQa278zldSO2UCTDdZXtBP9kAMIok3VpVb3kSWUnPjYlareFXy2
WcxI05OtKIEAlnSUZvy6292O0G5cp4UUIDIyWGkUQrAHm6HYGZN15qXTRaC5/t+fRgWq/oxqTWlf
XpxM5jXafITsHMt6wUKBMPD1AJiFKBVJT3zI6EO2OUeO4ekIRSd57wVQ53s6JdI2PVwegKUnY2kY
9zPbP7XWu8TAq8KdvtWypNtvoVYkQHrcKzUT1U/GCgiKxaPgbIOInYkpRV+O+n/5XgAol3w9VXnc
e5j7VcLdZ8OYcS0OAUsGzcRnsw038Y+CrP1BQr9a4qatl/VJe7OZioXg1RidFxH9OEL6T+mrmI0W
7qzzF1GEp/v2B188aT5hQIWTRkqjGPSnMXc3wi+gFkVjthD4Y7Slfkqmu+Uv2crPGfwSnM04Hv9h
YDidYYhca71/isJovNRFUrfC2PPYuUeuURYPepsry1NXg/3F0MLnPjII9N0uz5dLfyCM5nhc2YA6
WCDE9ijKaLlHqXS15NWmSF/9FORxfyB7Jxl7082izdK/aZjW/tahab0u++okUyaSFO9jBktdw9dB
ypYBzFwmazrzfQWyLDwxebmfmiMsRzyIbydxKORxxiNLCvXIS2dES+XhI6u4Jax3icR8JkV8ae7z
o6nur3NDInThIBOqVwds9pZU8NfhUR5pzQuSaEvuXBhB45XRMmhTS6tIyIP/7b+gfr+8PHm0wz/3
grBUwETT2Lr6EY2Mmy4udZ9wr3tVlhjKDYk6oNe6aYznqjSUE2uOT5nQx0da5aMTP8f79sLMMJgp
wqXCy7DVoo9TgBhMrq9CaO7BUrd0jlRm8GiNss78RRo9Tmr3AL4G+mTv1zqWJ41HZLAc9YYZ7w9T
cNIVMkKL58j8BLdM8cx/TFNxxCOfIxwMuOX++/5hycgdeaH29f2Bu5Cn9Q/Sym3aXyak/eBFAvIa
fPBPt7sYWLM+tH4CNz66VvLgvhcE+RJ6BrehRpvzHby3rdjZiQWXIzHUqbwMdlagQq+vMFf83n+m
cvzthe964BIcTFyXIjvwj51IETlg879wHoLUbbuP84Ja16duUX5HItIUUYOF0/iAvcw7Rm2YEDVy
1m0yjdJkgjzLruoaJZeCUjmCX7DFt4yVCRhkNrs/CjOfHdvhoXz7VTe/f36iIXpQ+1XrOmIL35Y2
Qwyw802U/tdghQZl8VojLLfvxVB39h27e4JsOUPBilr3WpenbD7bQ1mWurV52JwkInNMl2IX+xPB
uhMyRN3tD+JIvJgjYTu8BQvE0psJgR/RkiJtkrRcN9fTcvIu0OZSGQr5FnRhMj4+5zLpmKT8Kjvq
P5awqRh929vZR8dnbKDHZE2s73brBJbUveqUR27xQNdowdpJGZ5O/F4tUwfvhRGc1Vz9abBdoamh
LxiTSmfGZs6KAWA2TbR1l6r3u004u5tDAqwHwqK1LzeETCYGrcgjPJalqNun2Hdk20otuwFUB/Fw
8x5vomlIByfwqAp9f1MNsg50cR0RtNYGyja908L8JersNXXfOSml9+HRgbodmiMkksYttxt9Yqrr
RtuGTolLUYP4DIRmsVSDVD94Il+Y8dq101P6Zlyt4W9tZcKI21JIObVcNQL6oJT+idTvqBAYpP2W
ANMncXgUIV3YJaaJHFVd1K+PJZfKFZtIaqMXdt+9bKvDKaXOh48Tkl+tGod899W6SyxEF4vHm3fJ
w4n4buE3v6DpIgVIR3ZJVLJ96u95rdcNtFnzgYji37Yvt5UIsGqEFZ3OVeioabD+Yn3Ht/Mse4fW
jBW43Y67VGZ2kQzXG/razREzBBXVSB8adWa0zykxuZzyrXK020Ylom4m9zfK2cSAn+/57iabBl2B
dL4LcOOUW9Wa0RGVSysX6OJJbcw8bkeo+IRo26Ydz+b5Bsz9/0N7GokuwoNnaPLxDN95JZ1t38MB
wxIdLCV8rVnSOeS0Bz4U6X15KqyxYG0du4XyLf+VIBLkT2nt+CqQ72cjhqueKg9c4mdk9Nv/KTih
pdOD8JpfalIQOuiF7IsnDYueB0JIiuNaXiSxS/lGUUuUzLMAB+qfp2oiKg2Mck24Za+I/Kby3IW0
PsAEm+ju3X1vDsU8ly+L1YyRDmAnjkYA33FX0ztnSUaiHLnXRnb6Np54Hfsp3J4eGAhc2ygVKCMB
HjAxOacFFa/jnshYe/AK/shVXITojycw0aBz+N2QLokGdQpwM4RQ1xQ2g+068Axnv6aP3t7Sjqk1
u0eYm3jDYmvUHrr8IshUgUkawxYRdz/XN5nT8Qa32n1e7nTIFOjr/GwBGDAB8hIh60D+z/UpLKVa
zZeF47gqyA98XXdpxUm8jaafeLztDXo9Fn4I/KIomJjjuQtFBrrzXkvROWbpVE4A+itKXJeQdgUq
WNq9ZUZEP24wvirs+S+aQSDF8DibVjMKjTVqqcg2ClgTji83XRee1c4fhQ2pW3XRlQCHCnD3g37A
3lZVtXqNceFTFXWoZiUnlhOdI/ebm4PBWX8t+t+eZomBCkzMOr063Yxuhf02tkO+b5TmGsP0uhQj
W5plx5Q9RB7Mu3XMIQ/dYmmSvbj3WVTnSGCHwR1e0+l5nxSlf9PD6J8nzKlrsoG5SmF9Bn0Y+Ep5
NAWxpwUCb9XCM/3fTM1hH9tCUVoCvKlGOAx+rA/sbdwqnHBS1lPKJ5RHk12fUZADahrTSoX1a5BT
PO4tfpp25iw8KTbhoQghdXdOwO2xndYgshZ+m9X/1eVW7kaWGY1smCCmPN3zTOt69WKKUM/IAFFT
ihYnC+u+KF3KZO7YnnZLwwrQ8kG5mVzHM5jdT50GKkHqogIRVOVIUpW0kldHR1+HO3imSj9vi1zc
NY2ItLWX/KMRKe1Ywk64BF5JgRxUwdKkfMfnRAFM0lLxtQJH32WIdTPQzqv4b86XxNmP9Sow6g1e
kCdxE90iZPqhDLFhzEkmJXAVkQ9d1VaME6o1nT7yszY/cfJb2ZUIV018hjtbZmXWrCcjTB3o5dZH
jZ+gDgNCVCnIv4pAk3dmM2/hcEf+5TYUchMPjZkHleRjFqETZTApDypUF+6TZSBY/z0SXJquZGbU
45Rj3kUOiOIaT4mi8K6Hka+GOrhLI7crmO4CnEbD5WrdlWJVdHQWO+HCInhS2IsqBSmIMIBVLSn6
YSgNB+/bgSbER2+opdN/ZYmgprSc/nnTN9Rs+xHzdEPVvvi1J1rMjsHuNEDp7m/UQlx25TbKYDnE
cu9wE4Q9iGUTAyuYm+JV67FMtarZeNQheohQG5X6/z4rgaFrJeFBmyOGgX7xIggCDuB4MfuhwlaC
QRRPz3FqmMSo+yNaEYjfqBOSpbLH2Okfl0c+FdG0HvNyHVIQdUY1d8Ss2/bICxlOYvOL/CNkkzdM
DRWKsJE7+WatvNOxPJrcXgcUKi7WSWP7V7eakIcrd4w3T0k1Slm2/gNTlVmKiGB1PLiEEE3NjMQP
pqPoa6H96FXw2M2GoY7Er297xDfGP98ZIZsj48FTsRaU27NkZgJ9w/Wso1fUTpC0/v46ldKG3LMM
Y2fPmU0tU5z58qgbLkS6Lfdijdfe7R1rQORRrtMzh/4AK/UaCFI5A6QRq2dKdapU4VaxV0MlaIhL
Kr2RLrhXUTD1Xmkoh8TVCQREPMbpiknPxkjY2szhkyiE02YUQ2W8pEhQ7CferMDxZbZ7djUCrmFf
kqT4twdh4Cd2mG3F7OIZK12BCi8l1WWaMv3MFJdXgV20Zb0k7+UXb+aP3cwhB2/THuBqFtYK3tb1
8DswuZwd5ec0Jj+bHXF/z58zzJUj8wLXxTSSzPjrNHDcyr/LFoRsyFwsrkBQZ7XPv8I9CCG8iACI
TXkklDq281vvJD0fdtN5vIUKGKkqT09eprY0sqfVjgtqCFffJmhEzCJtSLq3cGGDtSxYBe8JPZTc
OtjhyG0Hr1+2J25jf+Lx65TaZoeoBSQM2CimqUQMt9GXRtyZ0PX+IbCQH4UmXwUTjjfRykDxP3oU
RbVEgtOVw509+lfWUNNYY96FDxfnH71oGC32GWy8z2HZvwGNPV+vE6dKSRGGKR7hiohTXJ/GT4U4
GRL3BCm3Jbna2yj4dT4xz0mj2064wJM7C+zTV/WoCYhzEGIgjAIMRiAxzarVQoA7ODt8zBcfkGkt
AE8VMBxaGZOQby4RLurAnf1KjSKFgs/xSue4nomNAzZJbAYmNTC9BZiPAHFie+3jvsv+iGrFuxJP
B2AELojJVGW83dca23U9l18o6Aw9/91xv1ZyMvhETIoATjwWR1LiciVJRj9OYtpC/oMjju5KfjS0
YR2IwC27VF++/D/owLJLhvmCAmELF5TFtFTblMC8vkn6eYDtqXIIYN+5nzQgmqIJRMRszfCAJ7+v
8/BNoHpYVIKThDWzu8afsyA306N/BljfhLns1j/LZfRKJ4r/BH2pqdkOX6L9fU92OdyN1NZJLrsh
tMzHftg3KUtRMg4XX70ppFNOrsM+6U+AJbXDsDGZVzRZcrqYwByS6rNjR4mhNJp3k7Eaev42y/Uk
L2SlSWrdzf3qiNLJRYr8yva3DRAkQaEkal9XeehctEOj/aczm+43KvlPOQX3jFtzW05sTpwjcKxn
8XCACaNMNZgxu87FjV09FDZfTHLBsN4uUbjgR3ICNxUmschqBk9DEg19h17nKiGV69ZDG8XDFFq9
/L+i+Wty8LZAJk05Wy8odw6PG6lKb1lexVWvxOlWIDyG/XdGTJwNXEe+huELqcIhQzrBpJl+z5a1
gb8y9QhlMwFwf8bjmTee8tr95rifoHt6he8OBzbZb3SPpS4JM27+9nupilH0F8wrGiNIEFql40+k
KwVJbu9vg93u9zA4Pg/gtBooAzYNY4V3Q7GxeK6kmg3ub8yMaiAt15wIx9piSx7YFT8Neb8QUUCb
Xthgr8c8i8p9AIrxIgnWrUcBI8m8S0dbdDSRwdHmtTjRwPHONMvlGTjys3IwExadwztaNHEVpLEM
uXqlqzMBNkVei/vX31vAPGmlNTpbWgoJXQi1vKe+V+XGM0FdXTzIf6LOM29wRSLs3KPfc/IoS8PY
/2cLhsCSloZ8zG25XoGnZhZoGMzjb3Szc5ugVQ82pdAmbLWBuPFLUJyMpu6f4fhQ9HVHv3bNjLxv
5eulRBfM5hgTepwLS25ZeqtVcm0Rb0sY8Ir6GKItu7CkTQMCPzZBDHkcORV4GGXO5u4cnNpHRnAJ
iiZPB+gjiUUwlBi0z/GsqhLxg4xnulNksK4t09ftRfbl+Vfc1ojdJetMDsSmA7rsKFLyOIg9WuK9
BYMinRA80jdY+fvJs3Bhw9Mn+jwj5r6G95nyz6JpJfs8q3e5Egu5gYboQD80o5SV7CnSqlFh3u7R
FvQAQ3r08ykkH8kB93+UjNz2YiiAhN7BwW4lmkN2vHa8Sq4N6k/SVqhchUQC3TEtlrNarAvFPDK8
SWKb7f4MQ/o4O0H22ywi+oncAY30mQghyfXzwbZ/TZ54KdmkaHyYEU2MEHxGoDXyUei2+SBQsE3J
kR0V4F8leMvYqjEMIymEguHN1pj2VwpmdnrzOTkmt5iCovcXnTV6qAitfb+lVLjO+eNOFnLzqaU7
F1WuAyWhQBW+mLl3uDHKVm5fSOi+Km+WH5LJJ4eUQk91Lu86SiikfwW3leiQ7ZFWlICNa1G6NQN7
3GivGBx++oeFlz1jIz7Uuwj9+YjzcaI0FU6iZdaGF9zpsbSCB3En8VvwVtZ3tA7uIlNnWuIwtpbC
rBVMXAuaFyyzV6UqMp43FQ8vBMxRY/Baa0b8oqmw3gtNxy1eVSBJrK9XybWP/6KMdlS8SqmubWpi
aYfCzG6a/HQPg75hJdpvongS2/cJBp0z54vOTJG8sv0wnFjTN7m3faKgOWYnWmT7BTB5BxDlEBG3
RvHapN5qQI9KKwiSpcymxsV5bc4U+GwzgSIko8rj/UG+VdsKPBlW+RYv1SY2JXqHDdHYCtB7UF7S
bmmZgDEnPDg626wYaoUHi9V7rRqJAjfZAZDIP5p4vzxNfs8Deve1bRlp45bIG7jsv8MeOseEOL/S
AG6BSl4KKudC3k07WiuJ+NxkClvZPsQzbNgK3krYfARKJJMrJHpazZMz/XMzcCgiAXavX5iqfPF3
wk1enSkRSqNvOEiuPwmypS5JZt0odHlIwmhGoaOoq3cCGh7Gx1zrgtktLawxeli76x9w9z1VW3cw
WCyk78HEvX6ryN/C9aFwZeDFVY0IDb9XMabNJ++HKO/ZO7ZbFzeKs6ol0ZEGm6pf4Qo9zU4O2W9+
XF5ku4ZRrQiaN/Py7OcQcObnbV1WDqqZvDtqjQElyvuGh0qkgCHg87YcVydDbf31LfDfLhOR09cJ
H/Kh0+E9fZursEMZS7egroTN2hd9ghorWhBaCXLaA/y8R502m9oCZhlU2TsLYp75a+Ojba6kt0qR
ht8sc4aUOk17lZLZ+crz9MUkXCtPoHIFa4zH7jhuENR5YJzJKmxU0aq3v9JDR+qMN2uwOydBitwB
59ZXqVKtvofVeSkH5Qry4I/YCbGQmNW2PQMWSxooNCS7MWYyiEOP/7lnu5sF6b6hMJ+MYYyNwppc
/fvhm5ySJB/51ODR4S7qp50Jc1lU9Y9NQOK9tfpySwD5ry41baASDF7S+iS8d/2K5r2B7VH5ngUN
nY4Tbhjyig3SU7l3Up8OrgwlBTTcYI5pMmlR6ZTOWIAWQzi6VyDnavvNRaL/2iVBTkl8puydrgWV
PmdetG0Frm/QGuqLUdNvfsR84eYri58A1nfknFiEKlvKmMjYIG2bBnkNwvg287t3MoRmvQv8CRZz
/DTxQfVUYtUJ4LCC4aCz1jAGkS0/BjKVw1qCNhI4m6yPf8mLo+HTWU1ucXM6WMOuHGTSKataVH+O
Ii6N7vevLdDcv2crzEHc6HiZHXLyjA+7LyvMPfDyDxVJBz6oH+OMYK8ODGklzhMgHVKzoqv2w7ZD
zdR/lG0OOuvGiTzx5jYY1XUgrTxlM7i1lXOF7A3zTh8+F9hXnK94U9RCPWUCk/nBMWakf5ec4qvT
SiUw4PKVmRfLtscIaaE4XqMDAzkENdWezbiptgvRC25tASFXfg2boZUZLcoLey/dKUAriMW6mG1C
8J2JEAbp4+WKch1PhtXtz4xP0mRD+IJ/ZZNbtdsnF6hpNud+zW3WqNy0yWrHXnJk19G00fkr2w24
ITx0HrN3FfRM937mLQBc8WkCca1oOEGvnqkz9FiM/1GJQNwB+tmSVHT0ReMSdp2WRfo8SuxMGMf0
SqEyFK8j8kbpDCroLZ/Ppw9/6mzgLRZRITJ7xBp5MRL14Dit8ARW3cFnE7Q9izz5tk7oYe5Hj67N
SkLk4yl0boKwm2MLY1FQnpqE6QjXJnBMMJFdYejobgFsKfSVOuIyUQTyTUyzAKd6PZuwvcynntKZ
DT7OeEGw2S+faPtnpkDhFgC0BHkOUESG2qRg6y78nw9h7xgbLn3vDjn6YrgCv+JKexvY2HqtQ5YV
GoTnmLWp48xZCWu+KN4LHyK9QZhqWMTLllvgtcSIxu5DqvlYCcqwzZWUh3i2Z2VoZWuGZeaBfasB
TZzi80uXsjvE8nCg9xvcD80bDiq4tr/mv8LMGP+8NKKYbUQ95m3zTo7Z/hWy9CpSx4hDLgIb9moX
L28UBdjQj1MMQuSkXQ98uGjSRIjCZy+JjoArTR/lB28ULqilu8KqzHmkMUfYPiwhjtjpIkISv7hN
pg2eheL8oVVDEyzuR0B+vpd13bXtPvZHHfDFXzmyOwZGj7mgrYssQ/qsuz1u+L8qEgT/Oi2p/wv+
tgn7YLKlYR40u6k6UAyqcnnF/eFypngElbXfVqfW2zUliV0YD3ptNJeMFvuypIIREKxRSgEhOTVq
OeF3hdgqITPtX+OQQvJRI2VA0IykZVjUxj3pOOpLSmgKMsyPqc9HjyKWE6sfZDVVlUcEEskOHJ5T
zx1lEi+xFuddRPqiA3rPHLB9lnRz60OraVQMMrfd1ks4xJNZM9FyfAYyXih+e2mAv5HUABETeSkP
Byoc50YteYbUscyZX6snZFzHRFb6TivKOUOPuLPNGcQWQeRv3f7pwPtPt4bH2wz8MMJJ7FSc4gVo
FihpFER7KxrEf5u+ZJ17XCsGG/kzcYd9ESzHUB8UZM3cmvu6jBRcfN1izf4pHXJFeRO9iL20ufuC
HsaRyvTkdoug2AnjTzEDPK/yQZT8gYDItjmAbpg7oVMSVgrtj+vpl7M9qvmAahs0rZPHWifukYgK
OsrL2U6n18JnoRchTqz3QRrXOwIeG70fojwmCmB3npTeIwXOw6feoPcIxT/kT5ZaeJJUpgTaonl6
hO83cPrAVWoZyywIO/vHBzdoaj4PqhKvcv6PMG7G6Hrr2VZs6Lnutpp75ODpQQyxdPuxYivY5/gi
BTrTiusCYZhSL9qrChI4c148K0C0LRO10aWl1rl0ftUBs92cEl1afJ6zwidtxhnbZaKQWRqccOI1
up4K6XUCzuCPlFpRUo0q33n6QFILO92qTiscSydD512KWU8kqZku1kcokTYnN/sXn8VJSDJes4E9
sJanGzM46UT1rL1S9PI92t4vYIdaDIKmpdPW50gPIHDWe8FCd3tUvMPrPhweDNrCGDesIVZ00snX
ZlUcKIVXtr6XgZPqEzjFi5eJJ6EV/ISj2fVjXsqqEi0WpkHfYvOYQSD7tDqakwkpUVQgivh8eC52
5wHcWTvYOnXceTfCjQDXKSKPj8Cg/AOAibBFielJU5h//sbb4uD4wOKXQD2FN0heFJF7oEht/9Sz
leGrYgPtxb86Rt/uFl4oEt4R6byBjVQBm+EgAcm5V6r+7fLXLyL0God/ddqrAhHlSOQOinF1gHqI
J6PmhOKGVVqhdxjJRLh5Wfe+2AWnsF6Q47tuowZPq+oqdS1oaKyJOsbKZFaPzLEHQv8UMscvj4/w
KRb59bvypKKKqoBhJva4eR0bPTLHyxMWN5s/50hFT+NYGdDctd5zadGGxrJmbJr9NugbDZYohvF4
hcdvm92ijGdm/B6PG1n2+cRKzzPhZymWnMCTOp3kEfPrZFLVwsdzsiwlNJA3/6PTz3j9LMwRQmPn
nL4kQ6WkJI6IdZKnOmrZl/rQFFMU2rILdsj4TF3HgkVx12bBLIt1qBCbjP/L3vKg0dakOrlc90Jq
vCudQscZfh9WnyGXGpzXMnC2YwH4ya6uYe6UnvrFj/XUFGi/uCHfanxPdhgv4w76plwKPWoB6zYV
6vGeEyMeT/U+DAfELmdxVleS+HYnBn6HZ2hwF25MYodi/9ZaKbUenm80rdFqtGJ2IhW0gJcF7v0o
y54xg/2ntqdPyqA+AhJr1CEI0TRNM8IjXjqJfRmTLwzxeNf1QDrJQfrZzrFIel8POyMDKsPi5HX+
R2cVRkIA9gjg4jh7X+A0djgo0Q3/ZVcB8l1bP2UKMxz++VSOQ56d6wyeNiBGBbn4yxdFB8mQm55X
+xs2CREBwPI2PTjx1wITrgIGcixZ/QeZayhY3LO1QD0PNU3srsfSFHUCIixJyHnKxMk1HnT2tA3U
TLiKwAz83DaheGnyDnnZP9gedEbGdMDXGVjv42qVFkJ7/qszbtalZpThLb+4FnUJ+68wbMrK+4it
AtBysW4Ubr0+Q3w+o78ACOh/0y10EZ4N0N6XOLsc01u7AqX/P31szjspp7Cl8rWz9uohYQLaKRYS
+tJiNDoH7KOtB43pcgxUhSNoSxujT4/i647NbrT7vQw5x9f2b6auFNuxX9GzPBA5e3jG8aLX2Fzk
PHYN6Oy6uBGDpVR8YH0FNMbZ7FcHrtiOFW+E499iC4byRqsTlwcVV5mXN4z6MqVoB9v1Pg8Y4HEu
qwGMI/tSzGElYZa7Px95gC0SRoSgsak9v7p5iZi5x/+5JS+fD/gj++iLPoFNcWUOOj32MyJCNFQr
Q15y1myt5MbROyTd3pkIyFK+NC4hm1hx7fwjTlBW40q4qg/AWKKWTFIrCqhZ0rsLpGgmcd3MyPHC
Qi+pdaAxSE/bzxHz9P20riLmxUy2vVucPChKQIvrlTQfOb3wD5TeNyQLJH/61//x4u+IcsbP8nFL
wF7cPEtb4a1pl2RuUmmdD9fVOjoecly8MpQdM8+izokvGCljir9deg4cN+eP6oly1/4klzA5NpN3
6Fi/4meER2f1E9yorSHvs56zA7E6JCqCQlZV7OEjV/UbfOiIu79DJ+pU0V1hI9EUpDNyKv5sUH5E
ZRW6b+QQX2Q9kjp3OuzYt0DX8JxAazupXIY2BNVjiLAVM0PXOmBri37uJJNvjdcrFAnQRJJVDK/K
aJNSbLQ6z8obqFcZeUJ2aYqmWpBP4r/CSwgxjiIPLYkgC80W18YWseG67qIgxic9rwpdXiLg2vtW
Lx086QvD474n/o2NgNaozf0KbBZtrrj+ER4hSaaNkGQ1la8xrom0gki8tMpmbXHU98VJQ2J5/SwV
pAiDzqDTeNye77m6AQ4bXMmYjdFKrJ7nHI1+3BY7ysEF9X8BlWB3zYW26WkVZ0tMe2diXXkFzhto
vo0UY3fGyTlFNFvBozDtzLUP3Qb4Vy3maGKHE52VVXWPSLJbS+CQX1VgGlOyA15zGtSqEDGQ/x2f
/jK7RG6+8E3InjTVAKgL8bbi4+HCoaDyUOsYrdtgAjXh1AwY7u2R9+fMoCSHLDP1X0TvWi0kgaUj
oCFai40dGPKijGgBb5xKPCrHPlTqJTrj7ZGfUTzLhBk3eRYF55AgXlZhcXkxeKPFto5U4ayryVFY
Jt7zhqueUTODxQ6hsmLbA524/zoZRXg/TWk14/qNIgFg2ZOhMD/VkkNP0rYUq0r9pEOpunRx6OHK
UfE8Mvq5iyuJ1YXDek/QUicdoZcwp7e9vkBAh05+uzww372ROSfq6G2nHDBQC5i0P4Ppg46XPsRQ
kSPv2OPxxUjOsDNjEIoKDvAq82W8f3bLf6kx0tTP/gOS/S6L3shjsnZs3g+v17mE1Go7ldlEBKx/
xG+nE2zmRZnQ0OOAgHCzandvLYJV76cJAgRaqZc52scMeYtiw6Vwq/DhIdq/sbO9F7sSpCfCvfK8
XHfmlcIxgd92QAz/fpmCi0icf2N9NOImdEi6mP17hi5RQDTh03JZ5me8mM9XvHcK5Ekf7tu5jI98
vWehtN5hrgx4+poUUA+U3vR802Sf4HsJCfvxh0b5C96/9REY+zUfJC+k4Ux3OynM/L7AHutm28qR
pcmwN/n/aTuUV2u1EYNijO4c40j9Z5xMHbk2/4JQfS1DPXl4mCSyDWcrN7t/Fl5bcAqpr/ame48E
zeFSEp4pQtzcnhk7kpydBklVehY2w0yFMQFzuVe6oxAOAuuZX2lcKbunUR7a0OptDqbnsyJj1te0
X9FoN60rRF5it083tvlcJyH+11Hlqhw839KZm2DD5o686ntIARdkqHGXXpEJPZSu9ZaL+Mp3BjQe
cXRUVMAUrqSHYXK//XAHaLbtlf4e3z7yAJo9xyzFDNu8aDRAtdDWtz99e4bTdeElHSJZjVjnJbwU
gWa4VBf8NBxOYgcn9SvaWXS6HcyilHaQO0oRJyIo2vsJcriOyZPJ9Zpo6hT6Rc8nI93hHZvXyz/H
fwPlHdPruMtaoV+ybcG55LP5Tf1tcDhl3PumiUv4+X46MooD1lFf1XhIkAjObe8o0gMD29QCAYQg
i4B9I8f1rZMmVPhp92AeFcOpPIJLW2HEHUs0TYJ0i1gX9oSfhpwj3ps5SyfdOdI8AYXv5P72TK1G
5MfNo1LhADoIxHPg74Yszy0RHkC+m+nmMcogtpMlwNSugj18CVFn/Gc4aShP8fiJNNxyrnmkIlcp
t3XsqnPAFs7jcCXHd/ef8QxVqRKz25cZmhziephHMfM60MXHLfhk9/JKxWsmanFy7tm1ZbmNPRYF
k8EPG9Ayyf4xfg73hpGj9CNjRUt9jv1JcLQeskqy/vHsxXOhV2RUPO94fE5IO9YJxPt848gvnt5m
eySJT1t1u6qrlBTfJcNPJQTMomtBTFoTJT6qhlr1KT9D4FAFqu5diROosA0ztBWCZTV5i2vHHQyk
OtDkMDamHuU3gQ7xheP4JLFBEQeyW0dRm1k1dkSgMsG6UEEHUYFlUAuQjo1F1Qtiu90GJoqCeimY
wMk6Kb1y3nfFvg3CVaGyhpRXXw0lwxDhZxwDQijHlCHrwHg4nCh2ky7ritApsZ31ZrkKXsY1zDi+
+FZTdSBPIPkbRtVyk7dY3ePpum9QYj0qOS2R3epi8NFgmTJS8pbwt1WrhBuoSLk3d35d87MaFJGg
qLr6jicx/Jl/3E7XDCbvW7P26uyUvEfAvWSUpfrRcGgrMO9QvgNtcGUohBqoV8qwO06qC9hJA/T+
F8aIlnYUrhKhBPhYnJAp0hzdM/vw6+pIzXQ4iwvFt3vFbXYbSJpnq2lSk9GKw83Q1yrT2tZRG7nI
iAWKDkkjvW1TC4lYYyI5oxKpM1HeviM9jaUmQlJ3WFV+NwXwDrT3aRii+C463KQ0hTidQpefIv6d
vCu47OgBImc4dpIrwNJhZlwrfQ40xNfrEDOtgwCmrBybIa/IegMzR7EYCthjyLOIpVHir1Fg0qZ5
Phpqf8pXphlXeI1du2CfefDurk8HpBM9B0QxrHfk36u/HPpQadmIBltZu7C5tdEs844XcVPWlDZY
N3yxCbUfWuCaT2mE7sXdfMdj8nlSqDQTdt1YDGo6VdnpQKBML0HUEiKaq3BhP4yKOPn16MVlM4yu
fU/VdE5SbsDWGxjO8w7zojwpOUvvfI6WAOKPnUSl3SFCLMYzPB/5e1SUAgX/l55VGhQ8RWogvYwW
J0VF3UvcyRAI5O9L89yqoH3WtiBtQ2EtTG6PPEU489/QK+IWYoyfFKX91REA/CQw6a58kil8JLrb
ut3kWPdUrPfEalpla57NNj4fy48iUD+mBfJjd3j5drS6AiPDfN4jGzpP26jcMrPrysCnkJ5wH5uw
4kSIhoSoM4Py2QLzNzCVLolM76otEi/EjKVlNPspACGrIenpAPFPlC2a5h6QGzfwGRi6FzJxQolW
DwBtoglGIhLPxc/C4M+L4XNhFSsH++ee3QBvhNtcc1G54Nj42vm39kKVyiLgKZPtVomtU8d8c8YO
cIgtTs6pA4mPMZ30hRmFGDLDpGlfHR6KSJ0oCVC6v+UDHpnWcVUnmiN+RGtV+slkbY5R9rZwdOTh
TgO+sx4g80ii4//xkNoksc9aGmOnVqfex9UgM3Qm/I4TO6I3HBxSS+/E+h9mJmx4stBp0WirdYFk
wHxMNLgpwRJV1Ruj67PM7fHi/l+aM8d7/BBQOoabjUBiKN0gWs6YSt3cs9kQyPPxhvTzCJDLh5ln
2VVdAGB5mRddz3Tqy3h7jE8/nnKrEXhzIp9hvEZ6ge3ZLp/yoZO/jf84YyBeI6YqwWhc9gCdL6bX
QUtvqskCvcZSqZ44j9K+n2Cqr0pLu3xD2AdOJTqo0q/vyxWn3vPrEvQ0cDAenDen5y2ITGcV6yb/
GPbqTIAvibnkSFqwNuUs1IztLeHD+s1Usnk8RXE5HrBqbs7hvWM4tSaDE6TqQGZo2NWngsBQPTkj
+WOr8HoQpPfqfxB7EpLAp4jeqBgtNuaaF5Q2Av4geeta6ULbL0io+gUc/QP9dPfAYOshriOzDGeD
dHEC4OVgiSFdBGpvCNWOwtOiFGPzTlfVc61CNqrEHIbLK4vaHZz6X9wNKXMD7cDmskoFXAPgAdxt
GUboIbYgFIx0KmTX+VAEE0daa81syvQ540ODeOAdIWheQ1YGqHhWIkD0x4FqiKuYKKq8Lph3KuSo
WsNYJ6KYeQE8yzqOGmYKfbJitfFoTE3aMWV0uzIi7zqKHQOhOyiik5itZUcSzjL2lmmhebiIseBA
FjYmc12Jx08cJJnB/LVW8yI4rvH4kUuYY/EkN0gdfnFY0xEseM2CWz5Nxe8NrBaiixkTpiFtaTuA
Aky52ymR0q9+qmERcdC8yZ3nJICMJDLu+Phn1WKDEyxByae2Cozsrcct90mVVQdFEyVJApr43qsU
Z+djWDa0Z+8NbDNuAqdcMSgvDZXhlAy8nFcgWK8dplRwWxrTYML2safsy38/p+OXBqXVkYPOX4U2
2Ql54BLfsS/smyBHPbrhZqzWNJTBBJvkC15vltgclu5pEMazbrI0/tuHWI/HKrEaY0N1IwB6YLPq
AV9qbK1z9bvMEqCjHOVwiRv707r77aEsL8TlCKE3T4YWxmhvQpHjGBoQyA2kcoPV+H7SidNwf1Wf
mxP2lbw5GI+Yu05lRRknC0BNv61rf79UQ+//527CQeBDV3L31Z4HIflIYwiYW0jmN+fIJgQfdM1N
zVqXTfgpPNVjDszALb5+vejiUvT2qoM+KQ+HZVaxJTlYz3rHVFYtup2ZDGsdLq1hdpFdSIEftkic
x9XADjWFTXwm9rLphr76tsX79AHWWIUmuM3D86pEnPgiWu9m2CaG5vcK/B3iPeeE/hOAjApGHklj
gkb6DhcDjghgNSg2eetSI/hXNhM2N2LRGZ5iTYURXcCnNejpxgi3dLIaD9nQK5hB3hVST7cbtYbQ
EOmxtt/PQU0MzkmL/z0123Vx8RYHpQR3D7tkTJYGPX9TA1bEYS6FIj6kkmezgrBSpKpHhlH2idCu
pbSKOm63OyJXtTQSeY3WIQcix/aMTpSUjFkmKiifJ3ZSqi6/wqU7hVBNg2jzUSkgZaMuUkUE+YZ2
+nmVbc5P/4JGGuN02bb4EKHwf/eWij/HH/lAGUz0avVSi/hvGIgyG5YaMgRkVEnIJSBmniGmONAo
VChJ8EyZqy4TQgjTnnEq1B1tAV1vISGsU9VGtsb0tTymBaYFeykHMFBcy+baZTjM8hYryyey2bZ/
+9kKz597FJtaqL0T8a/yUw6QF8cyPxZQFQj+3gw38sI53RBw0zjvFtZCzUkIRD0I1HdOHQzNZeDg
BojPmEZtta0DBP0goS/2NBWt75NzDC0/PrjbwHpUcCAsxsoSB/v5cJA9aqSnyVjhey+WQDpBs3IJ
VLSjKJ1kSxBpdvkMZSKEbeeDN3pYuz+0+Obcc9gHhHn2m0A6l1pBbxJhQsoiFHLDb79ykB2HPn6a
0pLh5HBRPObFz9RBLgwkfpb9uy3jIfaLGLA+w00X2dMRr53T5Pwlyvvq7q6gJWeN7tEBwOhpgNio
R/f4tgcrqmWfMCg7ca9m+976ixXRJ5hPNDP6fOrITKw/898Uovb3wnoMZ7eOdzYdsv9PcQ/ihB4b
mhXtWRe6OtGivMI0oPTlODMEZMz4Go/1yQ89RM0jvihpFJ7AQIr3wQ/22jJcOMTU9055ycF3d51g
+YQ4RDUcCXwKP5bhbzGLgmjUMxkterkjApkVEVZ9CoJ4HPf0HNah+CYk4FzOuev8or+ACcXz0umr
a14ZzK3FKqjxbABBkF0LzFZaXghyr1MBTSrfmoc96S2FHg1g1CQ1qAhdhbjy/2zGPPU5O+3AXctP
MCYQHNOYl4771pVcB8IRbusk6k2JCo3io5P2OKhZtaSBDnA8uy3UOFaysPgW6ruR8O5vskZVi80r
3NB7wWrK4h0X29jf2DdAA3qhR17e3p2AoYFmBTUt6MmgrR4bxbQR4MjkWdVpMBLuwhGb3ba6Jz3F
hdnh+/tl6pDB/viw9Umua78TqkDe2KQxqwubrp4IU+8MwD47gr7N7RgZT41nohNBbYhDob5FEqBU
5+/l3O+sKJb+crC/pRS0RPy+j8HpWexfwCcKIGw1Z4nS1rYSYm6eI8yEXttwMLUFLsBRT0kQ/2+f
z9Rv0fg/YKu4nN9QF7aVHcW3kL3mIgWM5AaOTyErehalLLtWa6nDC3aOORgtXFvegVzu2ZGrJLPf
bJ7UI11xua2PoPDX2bqF3Qtk9W3nqOe7gaDA98poogHQJskvK7ae1R/rBMr31Pej5nkCUn1jg9vo
LkqPz/87rO6fwPMONw6LT/0PuZMb0Q6UTKbkAOlG20yEnb1YXETXDDvheXEa+H2SElf+z93t5qfi
/z4gOGNEcMf91E94Fas6nSQnxuSGNnAfOL8fPHpc6x6uMRyQ2KBhS079Axycs7xoItyhI/q6f4Y1
g/oMq7PvQ6DgJmLp1yNnaLkvIFGS2yBphlcfqVPw5pwFc3CynkGJ42OigTMBDLn2aYHFRkkO4bly
UichPu7dFw6U2z9obi2+fD/S1Qmp8fFU7VAPUMYqwJAfrtE9icHjrQxVgk/8pQKxjR35BRfZIxwG
l76Qa/DUYOeVR1xtrSr2raDBif6j2GmfSUoZqHEBulOC7d55IhotDGaOmJfkHRxOscUr9DYmgo8Y
JIx1JbDylVGYcMVhbyH3lru8Jply2/gw6/I2C5JY1hjBs+/ZBc8B6aVf8RuIvB6wO/7orZ8RXCmx
cNnnutuftLuqROxE9XacD5UcMNMJJ6bre8R/CwZXmrsggHHSxTa7ZepzKukWO3mpqFX4fN+tZvKl
TvcqTx7wu+6iuUJJTuIVuoN+KtXhf3x7UXCuOeq34kGdX+VWTvkius5yJkfracQ7jiKmDGkNspcY
G3B9gxqZ1YzvheZ82hkPcdewbw7lWrBHCb/dQrv3FJ1A0c7V1jBPQDEGcBdURXdVEshpXo/c7nlx
CzbBnmecrRQud3cwqkfdlYWUH0BwciTG7mOT91sghVL/qwKVViR3U+xrQvrGnaNzHK489TUptt0b
E18c+D8OtnwbsXihv1NF+ORRXNsNJfhvC92nElnPt/zoai/u1rU52ubMoFllurNXW5f1rTzKTy2l
1mpfzzPe65hIUg9D1VyxEwXEXnilNOXEbeD02VTCrvcL8hLE19NxrYTWtKgQn1JyGfTW0HcGSTlt
yVvKwQYb+VyE5bjQhJOPRZiZ3fSnNLvm7kcrhkX2TLmkC/yuO24c+G76iOh9ChqrR1GUIFZD0ntN
NPXg2rwQ6MYnWmLu8xqI0hZjbcgq/muhNkzSGJry4UqZbUd+PkmVxAYXPSUAK0qbD09CvcvupYKU
pQ5jY+3QmeifNQXpWspkKOULcyqbKuaqA6McD7LH+tdcJ5moZUBnGA6hDEbQeJNOn2QRdRIYe/M8
elzfxMcguZlvvyKRyZlMy/B4J7YKae45XnTn2+UsUIbtCbtlgsyp/DhU1Yqe5QTSZ+iiW86WCZz7
vcnK1xBd+JMRA2geoyg3wPjD8cytcu6QiP4IfgvXp2kUK6rKixAIeTqvTCUAHpz6kmxMWqasr0I7
fNR5zI4KKVY3kLDnYJDojTMS4MFopzJhDiscfB5qjP5MJDVEj+miC/vAA1vfX9A9hO4+N464u4/0
3uM8iIzCn8X20VuHWpPQu88dEZBnDrkX3DVJuW68bFDu5ScJcb4gWrDzZ8vaE9hDAzEtwitG7P/2
APLo5fWT6YXK8rYNr7rnP7t4wgKbIl6w56IF7Pfb3y5hFczq4JF7oZCt7outLyCwe2SvzG3/nnhz
zRaRgSl2GMtHmnV58qepGqELgTiEQ+yZHyQecgAte1DPSpI/h7W2v+nl4J1mI7zRbff7b45yyotg
USRzLfabfUtHjK7wqvW7T+wAX+k+53UGVI3NAL1eBxJgLnNK871r9GtcNifmWxLytTkzH7qQ80CD
Q7f1ykkEeF3wj7c1sdequ3iGslfiNwJKU9ByyQchr3CFw2occDMj6oLgBZjQMonArevJtrM24Wka
TBbNZqn9yH8NstGgcYAg/moMXJmrBKvqQc+gg3KObWFHXbse47Cg4rVuROTTv8kBhDHc6WbSy3CF
MxczRVPEg54byUoUd34eCH5CRou8w3fogeQC5rEWQvGk+hzgn3qxd/+Escn0I4S8lnNZ+/GDUGa1
rwoDYwgE8BFIIlGacJdVj7ljxwAWQRyo8IM9ofNZGCLkW3gv+a9kdDdTUA1lPc3clQ6YOAvjHzPv
mU6K/2HPKbqIBQxP3sf0XMdIn8saMrxLbI+o/72OtZWUzVM5TGMn7xJF+jVPVNeHi8WMl/ow423p
L5zu2FMfG4RHPztdAVfpB/XMPEfJIzT8FUmie4zJljpIiEIypEM9XAwNQoFvl/VfFGGV6GGv8jlB
XXHBesKC4Msqaw4LdBt6/vuIyH3eZfMVF2GsQjgF12QS5nnazbRL10z0XcPEB+cYkfpSO4qZqjab
SSWF/FJmjqZd1kPE5B818obIm7Jx+amRvfwU5BIk9bWnrO/pr7HNxoLOD08sfmrDbKHTRks7e/R0
MQ4kLcIDEIfFPyKysGEqSD9nE3+QRBZSijTpeW1pLKdAFugsHj9aR9p1o2Hs/UYJFF3u1puhRKJP
Y5qqoz+DZnKMUqxGf3d8M0jCkCSUQZGE2DW6M9HfmOqqt8le7FSrQXx80bOIlFaElN1JQMhouy4e
dVil2wezAQ+1
`protect end_protected
